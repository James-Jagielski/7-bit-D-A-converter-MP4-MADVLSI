magic
tech sky130A
timestamp 1699841102
<< error_p >>
rect 15 472 35 475
rect 15 -92 18 472
rect 32 -92 35 472
rect 15 -95 35 -92
rect 215 472 235 475
rect 215 -92 218 472
rect 232 -92 235 472
rect 215 -95 235 -92
rect 415 472 435 475
rect 415 -92 418 472
rect 432 -92 435 472
rect 415 -95 435 -92
rect 815 472 835 475
rect 815 -92 818 472
rect 832 -92 835 472
rect 815 -95 835 -92
rect 1015 472 1035 475
rect 1015 -92 1018 472
rect 1032 -92 1035 472
rect 1015 -95 1035 -92
rect 1215 472 1235 475
rect 1215 -92 1218 472
rect 1232 -92 1235 472
rect 1215 -95 1235 -92
rect 15 -223 35 -220
rect 15 -787 18 -223
rect 32 -787 35 -223
rect 15 -790 35 -787
rect 515 -223 535 -220
rect 515 -787 518 -223
rect 532 -787 535 -223
rect 515 -790 535 -787
rect 715 -223 735 -220
rect 715 -787 718 -223
rect 732 -787 735 -223
rect 715 -790 735 -787
rect 1215 -223 1235 -220
rect 1215 -787 1218 -223
rect 1232 -787 1235 -223
rect 1215 -790 1235 -787
rect 515 -918 535 -915
rect 515 -1482 518 -918
rect 532 -1482 535 -918
rect 515 -1485 535 -1482
rect 715 -918 735 -915
rect 715 -1482 718 -918
rect 732 -1482 735 -918
rect 715 -1485 735 -1482
<< nwell >>
rect -20 -130 1270 510
<< nmos >>
rect 50 -805 100 -205
rect 150 -805 200 -205
rect 250 -805 300 -205
rect 450 -805 500 -205
rect 550 -805 600 -205
rect 650 -805 700 -205
rect 750 -805 800 -205
rect 950 -805 1000 -205
rect 1050 -805 1100 -205
rect 1150 -805 1200 -205
rect 50 -1500 100 -900
rect 150 -1500 200 -900
rect 250 -1500 300 -900
rect 350 -1500 400 -900
rect 550 -1500 600 -900
rect 650 -1500 700 -900
rect 850 -1500 900 -900
rect 950 -1500 1000 -900
rect 1050 -1500 1100 -900
rect 1150 -1500 1200 -900
rect 50 -2195 100 -1595
rect 150 -2195 200 -1595
rect 250 -2195 300 -1595
rect 350 -2195 400 -1595
rect 550 -2195 600 -1595
rect 650 -2195 700 -1595
rect 850 -2195 900 -1595
rect 950 -2195 1000 -1595
rect 1050 -2195 1100 -1595
rect 1150 -2195 1200 -1595
<< pmos >>
rect 50 -110 100 490
rect 150 -110 200 490
rect 250 -110 300 490
rect 350 -110 400 490
rect 450 -110 500 490
rect 750 -110 800 490
rect 850 -110 900 490
rect 950 -110 1000 490
rect 1050 -110 1100 490
rect 1150 -110 1200 490
<< ndiff >>
rect 0 -220 50 -205
rect 0 -790 15 -220
rect 35 -790 50 -220
rect 0 -805 50 -790
rect 100 -220 150 -205
rect 100 -790 115 -220
rect 135 -790 150 -220
rect 100 -805 150 -790
rect 200 -220 250 -205
rect 200 -790 215 -220
rect 235 -790 250 -220
rect 200 -805 250 -790
rect 300 -220 350 -205
rect 300 -790 315 -220
rect 335 -790 350 -220
rect 300 -805 350 -790
rect 400 -220 450 -205
rect 400 -790 415 -220
rect 435 -790 450 -220
rect 400 -805 450 -790
rect 500 -220 550 -205
rect 500 -790 515 -220
rect 535 -790 550 -220
rect 500 -805 550 -790
rect 600 -220 650 -205
rect 600 -790 615 -220
rect 635 -790 650 -220
rect 600 -805 650 -790
rect 700 -220 750 -205
rect 700 -790 715 -220
rect 735 -790 750 -220
rect 700 -805 750 -790
rect 800 -220 850 -205
rect 800 -790 815 -220
rect 835 -790 850 -220
rect 800 -805 850 -790
rect 900 -220 950 -205
rect 900 -790 915 -220
rect 935 -790 950 -220
rect 900 -805 950 -790
rect 1000 -220 1050 -205
rect 1000 -790 1015 -220
rect 1035 -790 1050 -220
rect 1000 -805 1050 -790
rect 1100 -220 1150 -205
rect 1100 -790 1115 -220
rect 1135 -790 1150 -220
rect 1100 -805 1150 -790
rect 1200 -220 1250 -205
rect 1200 -790 1215 -220
rect 1235 -790 1250 -220
rect 1200 -805 1250 -790
rect 0 -915 50 -900
rect 0 -1485 15 -915
rect 35 -1485 50 -915
rect 0 -1500 50 -1485
rect 100 -915 150 -900
rect 100 -1485 115 -915
rect 135 -1485 150 -915
rect 100 -1500 150 -1485
rect 200 -915 250 -900
rect 200 -1485 215 -915
rect 235 -1485 250 -915
rect 200 -1500 250 -1485
rect 300 -915 350 -900
rect 300 -1485 315 -915
rect 335 -1485 350 -915
rect 300 -1500 350 -1485
rect 400 -915 450 -900
rect 400 -1485 415 -915
rect 435 -1485 450 -915
rect 400 -1500 450 -1485
rect 500 -915 550 -900
rect 500 -1485 515 -915
rect 535 -1485 550 -915
rect 500 -1500 550 -1485
rect 600 -915 650 -900
rect 600 -1485 615 -915
rect 635 -1485 650 -915
rect 600 -1500 650 -1485
rect 700 -915 750 -900
rect 700 -1485 715 -915
rect 735 -1485 750 -915
rect 700 -1500 750 -1485
rect 800 -915 850 -900
rect 800 -1485 815 -915
rect 835 -1485 850 -915
rect 800 -1500 850 -1485
rect 900 -915 950 -900
rect 900 -1485 915 -915
rect 935 -1485 950 -915
rect 900 -1500 950 -1485
rect 1000 -915 1050 -900
rect 1000 -1485 1015 -915
rect 1035 -1485 1050 -915
rect 1000 -1500 1050 -1485
rect 1100 -915 1150 -900
rect 1100 -1485 1115 -915
rect 1135 -1485 1150 -915
rect 1100 -1500 1150 -1485
rect 1200 -915 1250 -900
rect 1200 -1485 1215 -915
rect 1235 -1485 1250 -915
rect 1200 -1500 1250 -1485
rect 0 -1610 50 -1595
rect 0 -2180 15 -1610
rect 35 -2180 50 -1610
rect 0 -2195 50 -2180
rect 100 -1610 150 -1595
rect 100 -2180 115 -1610
rect 135 -2180 150 -1610
rect 100 -2195 150 -2180
rect 200 -1610 250 -1595
rect 200 -2180 215 -1610
rect 235 -2180 250 -1610
rect 200 -2195 250 -2180
rect 300 -1610 350 -1595
rect 300 -2180 315 -1610
rect 335 -2180 350 -1610
rect 300 -2195 350 -2180
rect 400 -1610 450 -1595
rect 400 -2180 415 -1610
rect 435 -2180 450 -1610
rect 400 -2195 450 -2180
rect 500 -1610 550 -1595
rect 500 -2180 515 -1610
rect 535 -2180 550 -1610
rect 500 -2195 550 -2180
rect 600 -1610 650 -1595
rect 600 -2180 615 -1610
rect 635 -2180 650 -1610
rect 600 -2195 650 -2180
rect 700 -1610 750 -1595
rect 700 -2180 715 -1610
rect 735 -2180 750 -1610
rect 700 -2195 750 -2180
rect 800 -1610 850 -1595
rect 800 -2180 815 -1610
rect 835 -2180 850 -1610
rect 800 -2195 850 -2180
rect 900 -1610 950 -1595
rect 900 -2180 915 -1610
rect 935 -2180 950 -1610
rect 900 -2195 950 -2180
rect 1000 -1610 1050 -1595
rect 1000 -2180 1015 -1610
rect 1035 -2180 1050 -1610
rect 1000 -2195 1050 -2180
rect 1100 -1610 1150 -1595
rect 1100 -2180 1115 -1610
rect 1135 -2180 1150 -1610
rect 1100 -2195 1150 -2180
rect 1200 -1610 1250 -1595
rect 1200 -2180 1215 -1610
rect 1235 -2180 1250 -1610
rect 1200 -2195 1250 -2180
<< pdiff >>
rect 0 475 50 490
rect 0 -95 15 475
rect 35 -95 50 475
rect 0 -110 50 -95
rect 100 475 150 490
rect 100 -95 115 475
rect 135 -95 150 475
rect 100 -110 150 -95
rect 200 475 250 490
rect 200 -95 215 475
rect 235 -95 250 475
rect 200 -110 250 -95
rect 300 475 350 490
rect 300 -95 315 475
rect 335 -95 350 475
rect 300 -110 350 -95
rect 400 475 450 490
rect 400 -95 415 475
rect 435 -95 450 475
rect 400 -110 450 -95
rect 500 475 550 490
rect 500 -95 515 475
rect 535 -95 550 475
rect 700 475 750 490
rect 500 -110 550 -95
rect 700 -95 715 475
rect 735 -95 750 475
rect 700 -110 750 -95
rect 800 475 850 490
rect 800 -95 815 475
rect 835 -95 850 475
rect 800 -110 850 -95
rect 900 475 950 490
rect 900 -95 915 475
rect 935 -95 950 475
rect 900 -110 950 -95
rect 1000 475 1050 490
rect 1000 -95 1015 475
rect 1035 -95 1050 475
rect 1000 -110 1050 -95
rect 1100 475 1150 490
rect 1100 -95 1115 475
rect 1135 -95 1150 475
rect 1100 -110 1150 -95
rect 1200 475 1250 490
rect 1200 -95 1215 475
rect 1235 -95 1250 475
rect 1200 -110 1250 -95
<< ndiffc >>
rect 15 -790 35 -220
rect 115 -790 135 -220
rect 215 -790 235 -220
rect 315 -790 335 -220
rect 415 -790 435 -220
rect 515 -790 535 -220
rect 615 -790 635 -220
rect 715 -790 735 -220
rect 815 -790 835 -220
rect 915 -790 935 -220
rect 1015 -790 1035 -220
rect 1115 -790 1135 -220
rect 1215 -790 1235 -220
rect 15 -1485 35 -915
rect 115 -1485 135 -915
rect 215 -1485 235 -915
rect 315 -1485 335 -915
rect 415 -1485 435 -915
rect 515 -1485 535 -915
rect 615 -1485 635 -915
rect 715 -1485 735 -915
rect 815 -1485 835 -915
rect 915 -1485 935 -915
rect 1015 -1485 1035 -915
rect 1115 -1485 1135 -915
rect 1215 -1485 1235 -915
rect 15 -2180 35 -1610
rect 115 -2180 135 -1610
rect 215 -2180 235 -1610
rect 315 -2180 335 -1610
rect 415 -2180 435 -1610
rect 515 -2180 535 -1610
rect 615 -2180 635 -1610
rect 715 -2180 735 -1610
rect 815 -2180 835 -1610
rect 915 -2180 935 -1610
rect 1015 -2180 1035 -1610
rect 1115 -2180 1135 -1610
rect 1215 -2180 1235 -1610
<< pdiffc >>
rect 15 -95 35 475
rect 115 -95 135 475
rect 215 -95 235 475
rect 315 -95 335 475
rect 415 -95 435 475
rect 515 -95 535 475
rect 715 -95 735 475
rect 815 -95 835 475
rect 915 -95 935 475
rect 1015 -95 1035 475
rect 1115 -95 1135 475
rect 1215 -95 1235 475
<< poly >>
rect 50 490 100 505
rect 150 490 200 505
rect 250 490 300 505
rect 350 490 400 505
rect 450 490 500 505
rect 750 490 800 505
rect 850 490 900 505
rect 950 490 1000 505
rect 1050 490 1100 505
rect 1150 490 1200 505
rect 645 -35 685 -25
rect 645 -55 655 -35
rect 675 -55 685 -35
rect 50 -125 100 -110
rect 150 -125 200 -110
rect 250 -125 300 -110
rect 350 -125 400 -110
rect 450 -125 500 -110
rect 150 -135 500 -125
rect 150 -155 470 -135
rect 490 -155 500 -135
rect 150 -165 500 -155
rect 645 -150 685 -55
rect 750 -125 800 -110
rect 850 -125 900 -110
rect 950 -125 1000 -110
rect 1050 -125 1100 -110
rect 1150 -125 1200 -110
rect 750 -135 1100 -125
rect 645 -160 700 -150
rect 645 -180 670 -160
rect 690 -180 700 -160
rect 750 -155 865 -135
rect 885 -155 1100 -135
rect 750 -165 1100 -155
rect 645 -190 700 -180
rect 50 -205 100 -190
rect 150 -205 200 -190
rect 250 -205 300 -190
rect 450 -205 500 -190
rect 550 -205 600 -190
rect 650 -205 700 -190
rect 750 -205 800 -190
rect 950 -205 1000 -190
rect 1050 -205 1100 -190
rect 1150 -205 1200 -190
rect 50 -820 100 -805
rect 150 -820 200 -805
rect 250 -820 300 -805
rect 150 -860 300 -820
rect 450 -820 500 -805
rect 550 -820 600 -805
rect 650 -820 700 -805
rect 750 -820 800 -805
rect 450 -830 800 -820
rect 450 -850 515 -830
rect 535 -850 800 -830
rect 450 -860 800 -850
rect 950 -820 1000 -805
rect 1050 -820 1100 -805
rect 1150 -820 1200 -805
rect 950 -860 1100 -820
rect 50 -900 100 -885
rect 150 -900 200 -885
rect 250 -900 300 -885
rect 350 -900 400 -885
rect 550 -900 600 -885
rect 650 -900 700 -885
rect 850 -900 900 -885
rect 950 -900 1000 -885
rect 1050 -900 1100 -885
rect 1150 -900 1200 -885
rect 50 -1515 100 -1500
rect 150 -1515 200 -1500
rect 250 -1515 300 -1500
rect 350 -1515 400 -1500
rect 550 -1515 600 -1500
rect 650 -1515 700 -1500
rect 850 -1515 900 -1500
rect 950 -1515 1000 -1500
rect 1050 -1515 1100 -1500
rect 1150 -1515 1200 -1500
rect 150 -1555 1100 -1515
rect 50 -1595 100 -1580
rect 150 -1595 200 -1580
rect 250 -1595 300 -1580
rect 350 -1595 400 -1580
rect 550 -1595 600 -1580
rect 650 -1595 700 -1580
rect 850 -1595 900 -1580
rect 950 -1595 1000 -1580
rect 1050 -1595 1100 -1580
rect 1150 -1595 1200 -1580
rect 50 -2210 100 -2195
rect 150 -2210 200 -2195
rect 250 -2210 300 -2195
rect 350 -2210 400 -2195
rect 550 -2210 600 -2195
rect 650 -2210 700 -2195
rect 850 -2210 900 -2195
rect 950 -2210 1000 -2195
rect 1050 -2210 1100 -2195
rect 1150 -2210 1200 -2195
rect 150 -2250 1100 -2210
<< polycont >>
rect 655 -55 675 -35
rect 470 -155 490 -135
rect 670 -180 690 -160
rect 865 -155 885 -135
rect 515 -850 535 -830
<< locali >>
rect 125 505 425 525
rect 125 485 145 505
rect 405 485 425 505
rect 5 475 45 485
rect 5 -95 15 475
rect 35 -95 45 475
rect 5 -105 45 -95
rect 105 475 145 485
rect 105 -95 115 475
rect 135 -95 145 475
rect 105 -105 145 -95
rect 205 475 245 485
rect 205 -95 215 475
rect 235 -95 245 475
rect 205 -105 245 -95
rect 305 475 345 485
rect 305 -95 315 475
rect 335 -85 345 475
rect 405 475 445 485
rect 335 -95 385 -85
rect 305 -105 385 -95
rect 405 -95 415 475
rect 435 -95 445 475
rect 405 -105 445 -95
rect 505 475 545 485
rect 505 -95 515 475
rect 535 -95 545 475
rect 665 -25 685 525
rect 725 505 1125 525
rect 725 485 745 505
rect 1105 485 1125 505
rect 645 -35 685 -25
rect 645 -55 655 -35
rect 675 -55 685 -35
rect 645 -65 685 -55
rect 705 475 745 485
rect 705 -85 715 475
rect 505 -105 545 -95
rect 615 -95 715 -85
rect 735 -95 745 475
rect 615 -105 745 -95
rect 805 475 845 485
rect 805 -95 815 475
rect 835 -95 845 475
rect 805 -105 845 -95
rect 905 475 945 485
rect 905 -95 915 475
rect 935 -95 945 475
rect 905 -105 945 -95
rect 1005 475 1045 485
rect 1005 -95 1015 475
rect 1035 -95 1045 475
rect 1005 -105 1045 -95
rect 1105 475 1145 485
rect 1105 -95 1115 475
rect 1135 -95 1145 475
rect 1105 -105 1145 -95
rect 1205 475 1245 485
rect 1205 -95 1215 475
rect 1235 -95 1245 475
rect 1205 -105 1245 -95
rect 125 -170 145 -105
rect 125 -190 325 -170
rect 125 -210 145 -190
rect 305 -210 325 -190
rect 365 -210 385 -105
rect 615 -125 635 -105
rect 460 -135 635 -125
rect 460 -155 470 -135
rect 490 -145 635 -135
rect 490 -155 500 -145
rect 460 -165 500 -155
rect 615 -210 635 -145
rect 855 -135 895 -125
rect 660 -160 700 -150
rect 660 -180 670 -160
rect 690 -170 700 -160
rect 855 -155 865 -135
rect 885 -155 895 -135
rect 855 -165 895 -155
rect 690 -180 825 -170
rect 660 -190 825 -180
rect 805 -210 825 -190
rect 5 -220 45 -210
rect 5 -790 15 -220
rect 35 -790 45 -220
rect 5 -800 45 -790
rect 105 -220 145 -210
rect 105 -790 115 -220
rect 135 -790 145 -220
rect 105 -800 145 -790
rect 205 -220 245 -210
rect 205 -790 215 -220
rect 235 -790 245 -220
rect 205 -800 245 -790
rect 305 -220 345 -210
rect 305 -790 315 -220
rect 335 -790 345 -220
rect 365 -220 445 -210
rect 365 -230 415 -220
rect 305 -800 345 -790
rect 405 -790 415 -230
rect 435 -790 445 -220
rect 405 -800 445 -790
rect 505 -220 545 -210
rect 505 -790 515 -220
rect 535 -790 545 -220
rect 505 -800 545 -790
rect 605 -220 645 -210
rect 605 -790 615 -220
rect 635 -790 645 -220
rect 605 -800 645 -790
rect 705 -220 745 -210
rect 705 -790 715 -220
rect 735 -790 745 -220
rect 705 -800 745 -790
rect 805 -220 845 -210
rect 805 -790 815 -220
rect 835 -790 845 -220
rect 805 -800 845 -790
rect 15 -905 35 -800
rect 125 -905 145 -800
rect 215 -905 235 -800
rect 305 -865 325 -800
rect 425 -820 445 -800
rect 425 -830 545 -820
rect 865 -825 885 -165
rect 925 -190 1125 -170
rect 925 -210 945 -190
rect 1105 -210 1125 -190
rect 905 -220 945 -210
rect 905 -790 915 -220
rect 935 -790 945 -220
rect 905 -800 945 -790
rect 1005 -220 1045 -210
rect 1005 -790 1015 -220
rect 1035 -790 1045 -220
rect 1005 -800 1045 -790
rect 1105 -220 1145 -210
rect 1105 -790 1115 -220
rect 1135 -790 1145 -220
rect 1105 -800 1145 -790
rect 1205 -220 1245 -210
rect 1205 -790 1215 -220
rect 1235 -790 1245 -220
rect 1205 -800 1245 -790
rect 425 -840 515 -830
rect 505 -850 515 -840
rect 535 -850 545 -830
rect 505 -860 545 -850
rect 625 -845 885 -825
rect 305 -885 485 -865
rect 305 -905 325 -885
rect 5 -915 45 -905
rect 5 -1485 15 -915
rect 35 -1485 45 -915
rect 5 -1495 45 -1485
rect 105 -915 145 -905
rect 105 -1485 115 -915
rect 135 -1485 145 -915
rect 105 -1495 145 -1485
rect 205 -915 245 -905
rect 205 -1485 215 -915
rect 235 -1485 245 -915
rect 205 -1495 245 -1485
rect 305 -915 345 -905
rect 305 -1485 315 -915
rect 335 -1485 345 -915
rect 305 -1495 345 -1485
rect 405 -915 445 -905
rect 405 -1485 415 -915
rect 435 -1485 445 -915
rect 405 -1495 445 -1485
rect 15 -1600 35 -1495
rect 125 -1600 145 -1495
rect 215 -1600 235 -1495
rect 305 -1600 325 -1495
rect 425 -1600 445 -1495
rect 465 -1515 485 -885
rect 625 -905 645 -845
rect 925 -865 945 -800
rect 765 -885 945 -865
rect 505 -915 545 -905
rect 505 -1485 515 -915
rect 535 -1485 545 -915
rect 505 -1495 545 -1485
rect 605 -915 645 -905
rect 605 -1485 615 -915
rect 635 -1485 645 -915
rect 605 -1495 645 -1485
rect 705 -915 745 -905
rect 705 -1485 715 -915
rect 735 -1485 745 -915
rect 705 -1495 745 -1485
rect 765 -1515 785 -885
rect 925 -905 945 -885
rect 1015 -905 1035 -800
rect 1105 -905 1125 -800
rect 1215 -905 1235 -800
rect 465 -1535 785 -1515
rect 805 -915 845 -905
rect 805 -1485 815 -915
rect 835 -1485 845 -915
rect 805 -1495 845 -1485
rect 905 -915 945 -905
rect 905 -1485 915 -915
rect 935 -1485 945 -915
rect 905 -1495 945 -1485
rect 1005 -915 1045 -905
rect 1005 -1485 1015 -915
rect 1035 -1485 1045 -915
rect 1005 -1495 1045 -1485
rect 1105 -915 1145 -905
rect 1105 -1485 1115 -915
rect 1135 -1485 1145 -915
rect 1105 -1495 1145 -1485
rect 1205 -915 1245 -905
rect 1205 -1485 1215 -915
rect 1235 -1485 1245 -915
rect 1205 -1495 1245 -1485
rect 615 -1600 635 -1535
rect 805 -1600 825 -1495
rect 925 -1600 945 -1495
rect 1015 -1600 1035 -1495
rect 1105 -1600 1125 -1495
rect 1215 -1600 1235 -1495
rect 5 -1610 45 -1600
rect 5 -2180 15 -1610
rect 35 -2180 45 -1610
rect 5 -2190 45 -2180
rect 105 -1610 145 -1600
rect 105 -2180 115 -1610
rect 135 -2180 145 -1610
rect 105 -2190 145 -2180
rect 205 -1610 245 -1600
rect 205 -2180 215 -1610
rect 235 -2180 245 -1610
rect 205 -2190 245 -2180
rect 305 -1610 345 -1600
rect 305 -2180 315 -1610
rect 335 -2180 345 -1610
rect 305 -2190 345 -2180
rect 405 -1610 445 -1600
rect 405 -2180 415 -1610
rect 435 -2180 445 -1610
rect 405 -2190 445 -2180
rect 500 -1610 545 -1600
rect 500 -2180 515 -1610
rect 535 -2180 545 -1610
rect 500 -2190 545 -2180
rect 605 -1610 645 -1600
rect 605 -2180 615 -1610
rect 635 -2180 645 -1610
rect 605 -2190 645 -2180
rect 705 -1610 745 -1600
rect 705 -2180 715 -1610
rect 735 -2180 745 -1610
rect 705 -2190 745 -2180
rect 800 -1610 845 -1600
rect 800 -2180 815 -1610
rect 835 -2180 845 -1610
rect 800 -2190 845 -2180
rect 905 -1610 945 -1600
rect 905 -2180 915 -1610
rect 935 -2180 945 -1610
rect 905 -2190 945 -2180
rect 1005 -1610 1045 -1600
rect 1005 -2180 1015 -1610
rect 1035 -2180 1045 -1610
rect 1005 -2190 1045 -2180
rect 1105 -1610 1145 -1600
rect 1105 -2180 1115 -1610
rect 1135 -2180 1145 -1610
rect 1105 -2190 1145 -2180
rect 1205 -1610 1245 -1600
rect 1205 -2180 1215 -1610
rect 1235 -2180 1245 -1610
rect 1205 -2190 1245 -2180
rect 225 -2210 245 -2190
rect 415 -2210 435 -2190
rect 510 -2210 535 -2190
rect 715 -2210 735 -2190
rect 815 -2210 835 -2190
rect 1015 -2210 1035 -2190
rect 225 -2230 1035 -2210
<< viali >>
rect 15 -95 35 475
rect 215 -95 235 475
rect 415 -95 435 475
rect 815 -95 835 475
rect 1015 -95 1035 475
rect 1215 -95 1235 475
rect 15 -790 35 -220
rect 515 -790 535 -220
rect 715 -790 735 -220
rect 1215 -790 1235 -220
rect 515 -1485 535 -915
rect 715 -1485 735 -915
<< end >>

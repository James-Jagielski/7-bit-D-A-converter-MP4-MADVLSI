magic
tech sky130A
timestamp 1699851583
<< nmos >>
rect -5 0 45 600
rect 95 0 145 600
rect 195 0 245 600
rect 295 0 345 600
rect 395 0 445 600
rect 495 0 545 600
rect 695 0 745 600
rect 795 0 845 600
rect 895 0 945 600
rect 995 0 1045 600
rect 1095 0 1145 600
rect 1195 0 1245 600
rect 1395 0 1445 600
rect 1495 0 1545 600
rect 1595 0 1645 600
rect 1695 0 1745 600
rect 1795 0 1845 600
rect 1895 0 1945 600
rect 2095 0 2145 600
rect 2195 0 2245 600
rect 2295 0 2345 600
rect 2395 0 2445 600
rect 2495 0 2545 600
rect 2595 0 2645 600
rect 2795 0 2845 600
rect 2895 0 2945 600
rect 2995 0 3045 600
rect 3095 0 3145 600
rect 3195 0 3245 600
rect 3295 0 3345 600
rect 3495 0 3545 600
rect 3595 0 3645 600
rect 3695 0 3745 600
rect 3795 0 3845 600
rect 3895 0 3945 600
rect 3995 0 4045 600
rect 4195 0 4245 600
rect 4295 0 4345 600
rect 4395 0 4445 600
rect 4495 0 4545 600
rect 4595 0 4645 600
rect 4695 0 4745 600
rect 4795 0 4845 600
rect 4895 0 4945 600
rect -5 -695 45 -95
rect 95 -695 145 -95
rect 195 -695 245 -95
rect 295 -695 345 -95
rect 395 -695 445 -95
rect 495 -695 545 -95
rect 695 -695 745 -95
rect 795 -695 845 -95
rect 895 -695 945 -95
rect 995 -695 1045 -95
rect 1095 -695 1145 -95
rect 1195 -695 1245 -95
rect 1395 -695 1445 -95
rect 1495 -695 1545 -95
rect 1595 -695 1645 -95
rect 1695 -695 1745 -95
rect 1795 -695 1845 -95
rect 1895 -695 1945 -95
rect 2095 -695 2145 -95
rect 2195 -695 2245 -95
rect 2295 -695 2345 -95
rect 2395 -695 2445 -95
rect 2495 -695 2545 -95
rect 2595 -695 2645 -95
rect 2795 -695 2845 -95
rect 2895 -695 2945 -95
rect 2995 -695 3045 -95
rect 3095 -695 3145 -95
rect 3195 -695 3245 -95
rect 3295 -695 3345 -95
rect 3495 -695 3545 -95
rect 3595 -695 3645 -95
rect 3695 -695 3745 -95
rect 3795 -695 3845 -95
rect 3895 -695 3945 -95
rect 3995 -695 4045 -95
rect 4195 -695 4245 -95
rect 4295 -695 4345 -95
rect 4395 -695 4445 -95
rect 4495 -695 4545 -95
rect 4595 -695 4645 -95
rect 4695 -695 4745 -95
<< ndiff >>
rect -55 585 -5 600
rect -55 310 -40 585
rect -20 310 -5 585
rect -55 290 -5 310
rect -55 15 -40 290
rect -20 15 -5 290
rect -55 0 -5 15
rect 45 585 95 600
rect 45 310 60 585
rect 80 310 95 585
rect 45 290 95 310
rect 45 15 60 290
rect 80 15 95 290
rect 45 0 95 15
rect 145 585 195 600
rect 145 310 160 585
rect 180 310 195 585
rect 145 290 195 310
rect 145 15 160 290
rect 180 15 195 290
rect 145 0 195 15
rect 245 585 295 600
rect 245 310 260 585
rect 280 310 295 585
rect 245 290 295 310
rect 245 15 260 290
rect 280 15 295 290
rect 245 0 295 15
rect 345 585 395 600
rect 345 310 360 585
rect 380 310 395 585
rect 345 290 395 310
rect 345 15 360 290
rect 380 15 395 290
rect 345 0 395 15
rect 445 585 495 600
rect 445 310 460 585
rect 480 310 495 585
rect 445 290 495 310
rect 445 15 460 290
rect 480 15 495 290
rect 445 0 495 15
rect 545 585 595 600
rect 645 585 695 600
rect 545 310 560 585
rect 580 310 595 585
rect 645 310 660 585
rect 680 310 695 585
rect 545 290 595 310
rect 645 290 695 310
rect 545 15 560 290
rect 580 15 595 290
rect 645 15 660 290
rect 680 15 695 290
rect 545 0 595 15
rect 645 0 695 15
rect 745 585 795 600
rect 745 310 760 585
rect 780 310 795 585
rect 745 290 795 310
rect 745 15 760 290
rect 780 15 795 290
rect 745 0 795 15
rect 845 585 895 600
rect 845 310 860 585
rect 880 310 895 585
rect 845 290 895 310
rect 845 15 860 290
rect 880 15 895 290
rect 845 0 895 15
rect 945 585 995 600
rect 945 310 960 585
rect 980 310 995 585
rect 945 290 995 310
rect 945 15 960 290
rect 980 15 995 290
rect 945 0 995 15
rect 1045 585 1095 600
rect 1045 310 1060 585
rect 1080 310 1095 585
rect 1045 290 1095 310
rect 1045 15 1060 290
rect 1080 15 1095 290
rect 1045 0 1095 15
rect 1145 585 1195 600
rect 1145 310 1160 585
rect 1180 310 1195 585
rect 1145 290 1195 310
rect 1145 15 1160 290
rect 1180 15 1195 290
rect 1145 0 1195 15
rect 1245 585 1295 600
rect 1345 585 1395 600
rect 1245 310 1260 585
rect 1280 310 1295 585
rect 1345 310 1360 585
rect 1380 310 1395 585
rect 1245 290 1295 310
rect 1345 290 1395 310
rect 1245 15 1260 290
rect 1280 15 1295 290
rect 1345 15 1360 290
rect 1380 15 1395 290
rect 1245 0 1295 15
rect 1345 0 1395 15
rect 1445 585 1495 600
rect 1445 310 1460 585
rect 1480 310 1495 585
rect 1445 290 1495 310
rect 1445 15 1460 290
rect 1480 15 1495 290
rect 1445 0 1495 15
rect 1545 585 1595 600
rect 1545 310 1560 585
rect 1580 310 1595 585
rect 1545 290 1595 310
rect 1545 15 1560 290
rect 1580 15 1595 290
rect 1545 0 1595 15
rect 1645 585 1695 600
rect 1645 310 1660 585
rect 1680 310 1695 585
rect 1645 290 1695 310
rect 1645 15 1660 290
rect 1680 15 1695 290
rect 1645 0 1695 15
rect 1745 585 1795 600
rect 1745 310 1760 585
rect 1780 310 1795 585
rect 1745 290 1795 310
rect 1745 15 1760 290
rect 1780 15 1795 290
rect 1745 0 1795 15
rect 1845 585 1895 600
rect 1845 310 1860 585
rect 1880 310 1895 585
rect 1845 290 1895 310
rect 1845 15 1860 290
rect 1880 15 1895 290
rect 1845 0 1895 15
rect 1945 585 1995 600
rect 2045 585 2095 600
rect 1945 310 1960 585
rect 1980 310 1995 585
rect 2045 310 2060 585
rect 2080 310 2095 585
rect 1945 290 1995 310
rect 2045 290 2095 310
rect 1945 15 1960 290
rect 1980 15 1995 290
rect 2045 15 2060 290
rect 2080 15 2095 290
rect 1945 0 1995 15
rect 2045 0 2095 15
rect 2145 585 2195 600
rect 2145 310 2160 585
rect 2180 310 2195 585
rect 2145 290 2195 310
rect 2145 15 2160 290
rect 2180 15 2195 290
rect 2145 0 2195 15
rect 2245 585 2295 600
rect 2245 310 2260 585
rect 2280 310 2295 585
rect 2245 290 2295 310
rect 2245 15 2260 290
rect 2280 15 2295 290
rect 2245 0 2295 15
rect 2345 585 2395 600
rect 2345 310 2360 585
rect 2380 310 2395 585
rect 2345 290 2395 310
rect 2345 15 2360 290
rect 2380 15 2395 290
rect 2345 0 2395 15
rect 2445 585 2495 600
rect 2445 310 2460 585
rect 2480 310 2495 585
rect 2445 290 2495 310
rect 2445 15 2460 290
rect 2480 15 2495 290
rect 2445 0 2495 15
rect 2545 585 2595 600
rect 2545 310 2560 585
rect 2580 310 2595 585
rect 2545 290 2595 310
rect 2545 15 2560 290
rect 2580 15 2595 290
rect 2545 0 2595 15
rect 2645 585 2695 600
rect 2745 585 2795 600
rect 2645 310 2660 585
rect 2680 310 2695 585
rect 2745 310 2760 585
rect 2780 310 2795 585
rect 2645 290 2695 310
rect 2745 290 2795 310
rect 2645 15 2660 290
rect 2680 15 2695 290
rect 2745 15 2760 290
rect 2780 15 2795 290
rect 2645 0 2695 15
rect 2745 0 2795 15
rect 2845 585 2895 600
rect 2845 310 2860 585
rect 2880 310 2895 585
rect 2845 290 2895 310
rect 2845 15 2860 290
rect 2880 15 2895 290
rect 2845 0 2895 15
rect 2945 585 2995 600
rect 2945 310 2960 585
rect 2980 310 2995 585
rect 2945 290 2995 310
rect 2945 15 2960 290
rect 2980 15 2995 290
rect 2945 0 2995 15
rect 3045 585 3095 600
rect 3045 310 3060 585
rect 3080 310 3095 585
rect 3045 290 3095 310
rect 3045 15 3060 290
rect 3080 15 3095 290
rect 3045 0 3095 15
rect 3145 585 3195 600
rect 3145 310 3160 585
rect 3180 310 3195 585
rect 3145 290 3195 310
rect 3145 15 3160 290
rect 3180 15 3195 290
rect 3145 0 3195 15
rect 3245 585 3295 600
rect 3245 310 3260 585
rect 3280 310 3295 585
rect 3245 290 3295 310
rect 3245 15 3260 290
rect 3280 15 3295 290
rect 3245 0 3295 15
rect 3345 585 3395 600
rect 3445 585 3495 600
rect 3345 310 3360 585
rect 3380 310 3395 585
rect 3445 310 3460 585
rect 3480 310 3495 585
rect 3345 290 3395 310
rect 3445 290 3495 310
rect 3345 15 3360 290
rect 3380 15 3395 290
rect 3445 15 3460 290
rect 3480 15 3495 290
rect 3345 0 3395 15
rect 3445 0 3495 15
rect 3545 585 3595 600
rect 3545 310 3560 585
rect 3580 310 3595 585
rect 3545 290 3595 310
rect 3545 15 3560 290
rect 3580 15 3595 290
rect 3545 0 3595 15
rect 3645 585 3695 600
rect 3645 310 3660 585
rect 3680 310 3695 585
rect 3645 290 3695 310
rect 3645 15 3660 290
rect 3680 15 3695 290
rect 3645 0 3695 15
rect 3745 585 3795 600
rect 3745 310 3760 585
rect 3780 310 3795 585
rect 3745 290 3795 310
rect 3745 15 3760 290
rect 3780 15 3795 290
rect 3745 0 3795 15
rect 3845 585 3895 600
rect 3845 310 3860 585
rect 3880 310 3895 585
rect 3845 290 3895 310
rect 3845 15 3860 290
rect 3880 15 3895 290
rect 3845 0 3895 15
rect 3945 585 3995 600
rect 3945 310 3960 585
rect 3980 310 3995 585
rect 3945 290 3995 310
rect 3945 15 3960 290
rect 3980 15 3995 290
rect 3945 0 3995 15
rect 4045 585 4095 600
rect 4145 585 4195 600
rect 4045 310 4060 585
rect 4080 310 4095 585
rect 4145 310 4160 585
rect 4180 310 4195 585
rect 4045 290 4095 310
rect 4145 290 4195 310
rect 4045 15 4060 290
rect 4080 15 4095 290
rect 4145 15 4160 290
rect 4180 15 4195 290
rect 4045 0 4095 15
rect 4145 0 4195 15
rect 4245 585 4295 600
rect 4245 310 4260 585
rect 4280 310 4295 585
rect 4245 290 4295 310
rect 4245 15 4260 290
rect 4280 15 4295 290
rect 4245 0 4295 15
rect 4345 585 4395 600
rect 4345 310 4360 585
rect 4380 310 4395 585
rect 4345 290 4395 310
rect 4345 15 4360 290
rect 4380 15 4395 290
rect 4345 0 4395 15
rect 4445 585 4495 600
rect 4445 310 4460 585
rect 4480 310 4495 585
rect 4445 290 4495 310
rect 4445 15 4460 290
rect 4480 15 4495 290
rect 4445 0 4495 15
rect 4545 585 4595 600
rect 4545 310 4560 585
rect 4580 310 4595 585
rect 4545 290 4595 310
rect 4545 15 4560 290
rect 4580 15 4595 290
rect 4545 0 4595 15
rect 4645 585 4695 600
rect 4645 310 4660 585
rect 4680 310 4695 585
rect 4645 290 4695 310
rect 4645 15 4660 290
rect 4680 15 4695 290
rect 4645 0 4695 15
rect 4745 585 4795 600
rect 4745 310 4760 585
rect 4780 310 4795 585
rect 4745 290 4795 310
rect 4745 15 4760 290
rect 4780 15 4795 290
rect 4745 0 4795 15
rect 4845 585 4895 600
rect 4845 310 4860 585
rect 4880 310 4895 585
rect 4845 290 4895 310
rect 4845 15 4860 290
rect 4880 15 4895 290
rect 4845 0 4895 15
rect 4945 585 4995 600
rect 4945 310 4960 585
rect 4980 310 4995 585
rect 4945 290 4995 310
rect 4945 15 4960 290
rect 4980 15 4995 290
rect 4945 0 4995 15
rect -55 -110 -5 -95
rect -55 -385 -40 -110
rect -20 -385 -5 -110
rect -55 -405 -5 -385
rect -55 -680 -40 -405
rect -20 -680 -5 -405
rect -55 -695 -5 -680
rect 45 -110 95 -95
rect 45 -385 60 -110
rect 80 -385 95 -110
rect 45 -405 95 -385
rect 45 -680 60 -405
rect 80 -680 95 -405
rect 45 -695 95 -680
rect 145 -110 195 -95
rect 145 -385 160 -110
rect 180 -385 195 -110
rect 145 -405 195 -385
rect 145 -680 160 -405
rect 180 -680 195 -405
rect 145 -695 195 -680
rect 245 -110 295 -95
rect 245 -385 260 -110
rect 280 -385 295 -110
rect 245 -405 295 -385
rect 245 -680 260 -405
rect 280 -680 295 -405
rect 245 -695 295 -680
rect 345 -110 395 -95
rect 345 -385 360 -110
rect 380 -385 395 -110
rect 345 -405 395 -385
rect 345 -680 360 -405
rect 380 -680 395 -405
rect 345 -695 395 -680
rect 445 -110 495 -95
rect 445 -385 460 -110
rect 480 -385 495 -110
rect 445 -405 495 -385
rect 445 -680 460 -405
rect 480 -680 495 -405
rect 445 -695 495 -680
rect 545 -110 595 -95
rect 645 -110 695 -95
rect 545 -385 560 -110
rect 580 -385 595 -110
rect 645 -385 660 -110
rect 680 -385 695 -110
rect 545 -405 595 -385
rect 645 -405 695 -385
rect 545 -680 560 -405
rect 580 -680 595 -405
rect 645 -680 660 -405
rect 680 -680 695 -405
rect 545 -695 595 -680
rect 645 -695 695 -680
rect 745 -110 795 -95
rect 745 -385 760 -110
rect 780 -385 795 -110
rect 745 -405 795 -385
rect 745 -680 760 -405
rect 780 -680 795 -405
rect 745 -695 795 -680
rect 845 -110 895 -95
rect 845 -385 860 -110
rect 880 -385 895 -110
rect 845 -405 895 -385
rect 845 -680 860 -405
rect 880 -680 895 -405
rect 845 -695 895 -680
rect 945 -110 995 -95
rect 945 -385 960 -110
rect 980 -385 995 -110
rect 945 -405 995 -385
rect 945 -680 960 -405
rect 980 -680 995 -405
rect 945 -695 995 -680
rect 1045 -110 1095 -95
rect 1045 -385 1060 -110
rect 1080 -385 1095 -110
rect 1045 -405 1095 -385
rect 1045 -680 1060 -405
rect 1080 -680 1095 -405
rect 1045 -695 1095 -680
rect 1145 -110 1195 -95
rect 1145 -385 1160 -110
rect 1180 -385 1195 -110
rect 1145 -405 1195 -385
rect 1145 -680 1160 -405
rect 1180 -680 1195 -405
rect 1145 -695 1195 -680
rect 1245 -110 1295 -95
rect 1345 -110 1395 -95
rect 1245 -385 1260 -110
rect 1280 -385 1295 -110
rect 1345 -385 1360 -110
rect 1380 -385 1395 -110
rect 1245 -405 1295 -385
rect 1345 -405 1395 -385
rect 1245 -680 1260 -405
rect 1280 -680 1295 -405
rect 1345 -680 1360 -405
rect 1380 -680 1395 -405
rect 1245 -695 1295 -680
rect 1345 -695 1395 -680
rect 1445 -110 1495 -95
rect 1445 -385 1460 -110
rect 1480 -385 1495 -110
rect 1445 -405 1495 -385
rect 1445 -680 1460 -405
rect 1480 -680 1495 -405
rect 1445 -695 1495 -680
rect 1545 -110 1595 -95
rect 1545 -385 1560 -110
rect 1580 -385 1595 -110
rect 1545 -405 1595 -385
rect 1545 -680 1560 -405
rect 1580 -680 1595 -405
rect 1545 -695 1595 -680
rect 1645 -110 1695 -95
rect 1645 -385 1660 -110
rect 1680 -385 1695 -110
rect 1645 -405 1695 -385
rect 1645 -680 1660 -405
rect 1680 -680 1695 -405
rect 1645 -695 1695 -680
rect 1745 -110 1795 -95
rect 1745 -385 1760 -110
rect 1780 -385 1795 -110
rect 1745 -405 1795 -385
rect 1745 -680 1760 -405
rect 1780 -680 1795 -405
rect 1745 -695 1795 -680
rect 1845 -110 1895 -95
rect 1845 -385 1860 -110
rect 1880 -385 1895 -110
rect 1845 -405 1895 -385
rect 1845 -680 1860 -405
rect 1880 -680 1895 -405
rect 1845 -695 1895 -680
rect 1945 -110 1995 -95
rect 2045 -110 2095 -95
rect 1945 -385 1960 -110
rect 1980 -385 1995 -110
rect 2045 -385 2060 -110
rect 2080 -385 2095 -110
rect 1945 -405 1995 -385
rect 2045 -405 2095 -385
rect 1945 -680 1960 -405
rect 1980 -680 1995 -405
rect 2045 -680 2060 -405
rect 2080 -680 2095 -405
rect 1945 -695 1995 -680
rect 2045 -695 2095 -680
rect 2145 -110 2195 -95
rect 2145 -385 2160 -110
rect 2180 -385 2195 -110
rect 2145 -405 2195 -385
rect 2145 -680 2160 -405
rect 2180 -680 2195 -405
rect 2145 -695 2195 -680
rect 2245 -110 2295 -95
rect 2245 -385 2260 -110
rect 2280 -385 2295 -110
rect 2245 -405 2295 -385
rect 2245 -680 2260 -405
rect 2280 -680 2295 -405
rect 2245 -695 2295 -680
rect 2345 -110 2395 -95
rect 2345 -385 2360 -110
rect 2380 -385 2395 -110
rect 2345 -405 2395 -385
rect 2345 -680 2360 -405
rect 2380 -680 2395 -405
rect 2345 -695 2395 -680
rect 2445 -110 2495 -95
rect 2445 -385 2460 -110
rect 2480 -385 2495 -110
rect 2445 -405 2495 -385
rect 2445 -680 2460 -405
rect 2480 -680 2495 -405
rect 2445 -695 2495 -680
rect 2545 -110 2595 -95
rect 2545 -385 2560 -110
rect 2580 -385 2595 -110
rect 2545 -405 2595 -385
rect 2545 -680 2560 -405
rect 2580 -680 2595 -405
rect 2545 -695 2595 -680
rect 2645 -110 2695 -95
rect 2745 -110 2795 -95
rect 2645 -385 2660 -110
rect 2680 -385 2695 -110
rect 2745 -385 2760 -110
rect 2780 -385 2795 -110
rect 2645 -405 2695 -385
rect 2745 -405 2795 -385
rect 2645 -680 2660 -405
rect 2680 -680 2695 -405
rect 2745 -680 2760 -405
rect 2780 -680 2795 -405
rect 2645 -695 2695 -680
rect 2745 -695 2795 -680
rect 2845 -110 2895 -95
rect 2845 -385 2860 -110
rect 2880 -385 2895 -110
rect 2845 -405 2895 -385
rect 2845 -680 2860 -405
rect 2880 -680 2895 -405
rect 2845 -695 2895 -680
rect 2945 -110 2995 -95
rect 2945 -385 2960 -110
rect 2980 -385 2995 -110
rect 2945 -405 2995 -385
rect 2945 -680 2960 -405
rect 2980 -680 2995 -405
rect 2945 -695 2995 -680
rect 3045 -110 3095 -95
rect 3045 -385 3060 -110
rect 3080 -385 3095 -110
rect 3045 -405 3095 -385
rect 3045 -680 3060 -405
rect 3080 -680 3095 -405
rect 3045 -695 3095 -680
rect 3145 -110 3195 -95
rect 3145 -385 3160 -110
rect 3180 -385 3195 -110
rect 3145 -405 3195 -385
rect 3145 -680 3160 -405
rect 3180 -680 3195 -405
rect 3145 -695 3195 -680
rect 3245 -110 3295 -95
rect 3245 -385 3260 -110
rect 3280 -385 3295 -110
rect 3245 -405 3295 -385
rect 3245 -680 3260 -405
rect 3280 -680 3295 -405
rect 3245 -695 3295 -680
rect 3345 -110 3395 -95
rect 3445 -110 3495 -95
rect 3345 -385 3360 -110
rect 3380 -385 3395 -110
rect 3445 -385 3460 -110
rect 3480 -385 3495 -110
rect 3345 -405 3395 -385
rect 3445 -405 3495 -385
rect 3345 -680 3360 -405
rect 3380 -680 3395 -405
rect 3445 -680 3460 -405
rect 3480 -680 3495 -405
rect 3345 -695 3395 -680
rect 3445 -695 3495 -680
rect 3545 -110 3595 -95
rect 3545 -385 3560 -110
rect 3580 -385 3595 -110
rect 3545 -405 3595 -385
rect 3545 -680 3560 -405
rect 3580 -680 3595 -405
rect 3545 -695 3595 -680
rect 3645 -110 3695 -95
rect 3645 -385 3660 -110
rect 3680 -385 3695 -110
rect 3645 -405 3695 -385
rect 3645 -680 3660 -405
rect 3680 -680 3695 -405
rect 3645 -695 3695 -680
rect 3745 -110 3795 -95
rect 3745 -385 3760 -110
rect 3780 -385 3795 -110
rect 3745 -405 3795 -385
rect 3745 -680 3760 -405
rect 3780 -680 3795 -405
rect 3745 -695 3795 -680
rect 3845 -110 3895 -95
rect 3845 -385 3860 -110
rect 3880 -385 3895 -110
rect 3845 -405 3895 -385
rect 3845 -680 3860 -405
rect 3880 -680 3895 -405
rect 3845 -695 3895 -680
rect 3945 -110 3995 -95
rect 3945 -385 3960 -110
rect 3980 -385 3995 -110
rect 3945 -405 3995 -385
rect 3945 -680 3960 -405
rect 3980 -680 3995 -405
rect 3945 -695 3995 -680
rect 4045 -110 4095 -95
rect 4145 -110 4195 -95
rect 4045 -385 4060 -110
rect 4080 -385 4095 -110
rect 4145 -385 4160 -110
rect 4180 -385 4195 -110
rect 4045 -405 4095 -385
rect 4145 -405 4195 -385
rect 4045 -680 4060 -405
rect 4080 -680 4095 -405
rect 4145 -680 4160 -405
rect 4180 -680 4195 -405
rect 4045 -695 4095 -680
rect 4145 -695 4195 -680
rect 4245 -110 4295 -95
rect 4245 -385 4260 -110
rect 4280 -385 4295 -110
rect 4245 -405 4295 -385
rect 4245 -680 4260 -405
rect 4280 -680 4295 -405
rect 4245 -695 4295 -680
rect 4345 -110 4395 -95
rect 4345 -385 4360 -110
rect 4380 -385 4395 -110
rect 4345 -405 4395 -385
rect 4345 -680 4360 -405
rect 4380 -680 4395 -405
rect 4345 -695 4395 -680
rect 4445 -110 4495 -95
rect 4445 -385 4460 -110
rect 4480 -385 4495 -110
rect 4445 -405 4495 -385
rect 4445 -680 4460 -405
rect 4480 -680 4495 -405
rect 4445 -695 4495 -680
rect 4545 -110 4595 -95
rect 4545 -385 4560 -110
rect 4580 -385 4595 -110
rect 4545 -405 4595 -385
rect 4545 -680 4560 -405
rect 4580 -680 4595 -405
rect 4545 -695 4595 -680
rect 4645 -110 4695 -95
rect 4645 -385 4660 -110
rect 4680 -385 4695 -110
rect 4645 -405 4695 -385
rect 4645 -680 4660 -405
rect 4680 -680 4695 -405
rect 4645 -695 4695 -680
rect 4745 -110 4795 -95
rect 4745 -385 4760 -110
rect 4780 -385 4795 -110
rect 4745 -405 4795 -385
rect 4745 -680 4760 -405
rect 4780 -680 4795 -405
rect 4745 -695 4795 -680
<< ndiffc >>
rect -40 310 -20 585
rect -40 15 -20 290
rect 60 310 80 585
rect 60 15 80 290
rect 160 310 180 585
rect 160 15 180 290
rect 260 310 280 585
rect 260 15 280 290
rect 360 310 380 585
rect 360 15 380 290
rect 460 310 480 585
rect 460 15 480 290
rect 560 310 580 585
rect 660 310 680 585
rect 560 15 580 290
rect 660 15 680 290
rect 760 310 780 585
rect 760 15 780 290
rect 860 310 880 585
rect 860 15 880 290
rect 960 310 980 585
rect 960 15 980 290
rect 1060 310 1080 585
rect 1060 15 1080 290
rect 1160 310 1180 585
rect 1160 15 1180 290
rect 1260 310 1280 585
rect 1360 310 1380 585
rect 1260 15 1280 290
rect 1360 15 1380 290
rect 1460 310 1480 585
rect 1460 15 1480 290
rect 1560 310 1580 585
rect 1560 15 1580 290
rect 1660 310 1680 585
rect 1660 15 1680 290
rect 1760 310 1780 585
rect 1760 15 1780 290
rect 1860 310 1880 585
rect 1860 15 1880 290
rect 1960 310 1980 585
rect 2060 310 2080 585
rect 1960 15 1980 290
rect 2060 15 2080 290
rect 2160 310 2180 585
rect 2160 15 2180 290
rect 2260 310 2280 585
rect 2260 15 2280 290
rect 2360 310 2380 585
rect 2360 15 2380 290
rect 2460 310 2480 585
rect 2460 15 2480 290
rect 2560 310 2580 585
rect 2560 15 2580 290
rect 2660 310 2680 585
rect 2760 310 2780 585
rect 2660 15 2680 290
rect 2760 15 2780 290
rect 2860 310 2880 585
rect 2860 15 2880 290
rect 2960 310 2980 585
rect 2960 15 2980 290
rect 3060 310 3080 585
rect 3060 15 3080 290
rect 3160 310 3180 585
rect 3160 15 3180 290
rect 3260 310 3280 585
rect 3260 15 3280 290
rect 3360 310 3380 585
rect 3460 310 3480 585
rect 3360 15 3380 290
rect 3460 15 3480 290
rect 3560 310 3580 585
rect 3560 15 3580 290
rect 3660 310 3680 585
rect 3660 15 3680 290
rect 3760 310 3780 585
rect 3760 15 3780 290
rect 3860 310 3880 585
rect 3860 15 3880 290
rect 3960 310 3980 585
rect 3960 15 3980 290
rect 4060 310 4080 585
rect 4160 310 4180 585
rect 4060 15 4080 290
rect 4160 15 4180 290
rect 4260 310 4280 585
rect 4260 15 4280 290
rect 4360 310 4380 585
rect 4360 15 4380 290
rect 4460 310 4480 585
rect 4460 15 4480 290
rect 4560 310 4580 585
rect 4560 15 4580 290
rect 4660 310 4680 585
rect 4660 15 4680 290
rect 4760 310 4780 585
rect 4760 15 4780 290
rect 4860 310 4880 585
rect 4860 15 4880 290
rect 4960 310 4980 585
rect 4960 15 4980 290
rect -40 -385 -20 -110
rect -40 -680 -20 -405
rect 60 -385 80 -110
rect 60 -680 80 -405
rect 160 -385 180 -110
rect 160 -680 180 -405
rect 260 -385 280 -110
rect 260 -680 280 -405
rect 360 -385 380 -110
rect 360 -680 380 -405
rect 460 -385 480 -110
rect 460 -680 480 -405
rect 560 -385 580 -110
rect 660 -385 680 -110
rect 560 -680 580 -405
rect 660 -680 680 -405
rect 760 -385 780 -110
rect 760 -680 780 -405
rect 860 -385 880 -110
rect 860 -680 880 -405
rect 960 -385 980 -110
rect 960 -680 980 -405
rect 1060 -385 1080 -110
rect 1060 -680 1080 -405
rect 1160 -385 1180 -110
rect 1160 -680 1180 -405
rect 1260 -385 1280 -110
rect 1360 -385 1380 -110
rect 1260 -680 1280 -405
rect 1360 -680 1380 -405
rect 1460 -385 1480 -110
rect 1460 -680 1480 -405
rect 1560 -385 1580 -110
rect 1560 -680 1580 -405
rect 1660 -385 1680 -110
rect 1660 -680 1680 -405
rect 1760 -385 1780 -110
rect 1760 -680 1780 -405
rect 1860 -385 1880 -110
rect 1860 -680 1880 -405
rect 1960 -385 1980 -110
rect 2060 -385 2080 -110
rect 1960 -680 1980 -405
rect 2060 -680 2080 -405
rect 2160 -385 2180 -110
rect 2160 -680 2180 -405
rect 2260 -385 2280 -110
rect 2260 -680 2280 -405
rect 2360 -385 2380 -110
rect 2360 -680 2380 -405
rect 2460 -385 2480 -110
rect 2460 -680 2480 -405
rect 2560 -385 2580 -110
rect 2560 -680 2580 -405
rect 2660 -385 2680 -110
rect 2760 -385 2780 -110
rect 2660 -680 2680 -405
rect 2760 -680 2780 -405
rect 2860 -385 2880 -110
rect 2860 -680 2880 -405
rect 2960 -385 2980 -110
rect 2960 -680 2980 -405
rect 3060 -385 3080 -110
rect 3060 -680 3080 -405
rect 3160 -385 3180 -110
rect 3160 -680 3180 -405
rect 3260 -385 3280 -110
rect 3260 -680 3280 -405
rect 3360 -385 3380 -110
rect 3460 -385 3480 -110
rect 3360 -680 3380 -405
rect 3460 -680 3480 -405
rect 3560 -385 3580 -110
rect 3560 -680 3580 -405
rect 3660 -385 3680 -110
rect 3660 -680 3680 -405
rect 3760 -385 3780 -110
rect 3760 -680 3780 -405
rect 3860 -385 3880 -110
rect 3860 -680 3880 -405
rect 3960 -385 3980 -110
rect 3960 -680 3980 -405
rect 4060 -385 4080 -110
rect 4160 -385 4180 -110
rect 4060 -680 4080 -405
rect 4160 -680 4180 -405
rect 4260 -385 4280 -110
rect 4260 -680 4280 -405
rect 4360 -385 4380 -110
rect 4360 -680 4380 -405
rect 4460 -385 4480 -110
rect 4460 -680 4480 -405
rect 4560 -385 4580 -110
rect 4560 -680 4580 -405
rect 4660 -385 4680 -110
rect 4660 -680 4680 -405
rect 4760 -385 4780 -110
rect 4760 -680 4780 -405
<< psubdiff >>
rect -105 585 -55 600
rect -105 310 -90 585
rect -70 310 -55 585
rect -105 290 -55 310
rect -105 15 -90 290
rect -70 15 -55 290
rect -105 0 -55 15
rect 595 585 645 600
rect 595 310 610 585
rect 630 310 645 585
rect 595 290 645 310
rect 595 15 610 290
rect 630 15 645 290
rect 595 0 645 15
rect 1295 585 1345 600
rect 1295 310 1310 585
rect 1330 310 1345 585
rect 1295 290 1345 310
rect 1295 15 1310 290
rect 1330 15 1345 290
rect 1295 0 1345 15
rect 1995 585 2045 600
rect 1995 310 2010 585
rect 2030 310 2045 585
rect 1995 290 2045 310
rect 1995 15 2010 290
rect 2030 15 2045 290
rect 1995 0 2045 15
rect 2695 585 2745 600
rect 2695 310 2710 585
rect 2730 310 2745 585
rect 2695 290 2745 310
rect 2695 15 2710 290
rect 2730 15 2745 290
rect 2695 0 2745 15
rect 3395 585 3445 600
rect 3395 310 3410 585
rect 3430 310 3445 585
rect 3395 290 3445 310
rect 3395 15 3410 290
rect 3430 15 3445 290
rect 3395 0 3445 15
rect 4095 585 4145 600
rect 4095 310 4110 585
rect 4130 310 4145 585
rect 4095 290 4145 310
rect 4095 15 4110 290
rect 4130 15 4145 290
rect 4095 0 4145 15
rect -105 -110 -55 -95
rect -105 -385 -90 -110
rect -70 -385 -55 -110
rect -105 -405 -55 -385
rect -105 -680 -90 -405
rect -70 -680 -55 -405
rect -105 -695 -55 -680
rect 595 -110 645 -95
rect 595 -385 610 -110
rect 630 -385 645 -110
rect 595 -405 645 -385
rect 595 -680 610 -405
rect 630 -680 645 -405
rect 595 -695 645 -680
rect 1295 -110 1345 -95
rect 1295 -385 1310 -110
rect 1330 -385 1345 -110
rect 1295 -405 1345 -385
rect 1295 -680 1310 -405
rect 1330 -680 1345 -405
rect 1295 -695 1345 -680
rect 1995 -110 2045 -95
rect 1995 -385 2010 -110
rect 2030 -385 2045 -110
rect 1995 -405 2045 -385
rect 1995 -680 2010 -405
rect 2030 -680 2045 -405
rect 1995 -695 2045 -680
rect 2695 -110 2745 -95
rect 2695 -385 2710 -110
rect 2730 -385 2745 -110
rect 2695 -405 2745 -385
rect 2695 -680 2710 -405
rect 2730 -680 2745 -405
rect 2695 -695 2745 -680
rect 3395 -110 3445 -95
rect 3395 -385 3410 -110
rect 3430 -385 3445 -110
rect 3395 -405 3445 -385
rect 3395 -680 3410 -405
rect 3430 -680 3445 -405
rect 3395 -695 3445 -680
rect 4095 -110 4145 -95
rect 4095 -385 4110 -110
rect 4130 -385 4145 -110
rect 4095 -405 4145 -385
rect 4095 -680 4110 -405
rect 4130 -680 4145 -405
rect 4095 -695 4145 -680
<< psubdiffcont >>
rect -90 310 -70 585
rect -90 15 -70 290
rect 610 310 630 585
rect 610 15 630 290
rect 1310 310 1330 585
rect 1310 15 1330 290
rect 2010 310 2030 585
rect 2010 15 2030 290
rect 2710 310 2730 585
rect 2710 15 2730 290
rect 3410 310 3430 585
rect 3410 15 3430 290
rect 4110 310 4130 585
rect 4110 15 4130 290
rect -90 -385 -70 -110
rect -90 -680 -70 -405
rect 610 -385 630 -110
rect 610 -680 630 -405
rect 1310 -385 1330 -110
rect 1310 -680 1330 -405
rect 2010 -385 2030 -110
rect 2010 -680 2030 -405
rect 2710 -385 2730 -110
rect 2710 -680 2730 -405
rect 3410 -385 3430 -110
rect 3410 -680 3430 -405
rect 4110 -385 4130 -110
rect 4110 -680 4130 -405
<< poly >>
rect -165 640 145 655
rect 95 630 145 640
rect 395 640 845 655
rect 395 630 445 640
rect 95 615 445 630
rect 795 630 845 640
rect 1095 640 1545 655
rect 1095 630 1145 640
rect 795 615 1145 630
rect 1495 630 1545 640
rect 1795 640 2245 655
rect 1795 630 1845 640
rect 1495 615 1845 630
rect 2195 630 2245 640
rect 2495 640 2945 655
rect 2495 630 2545 640
rect 2195 615 2545 630
rect 2895 630 2945 640
rect 3195 640 3645 655
rect 3195 630 3245 640
rect 2895 615 3245 630
rect 3595 630 3645 640
rect 3895 640 4445 655
rect 3895 630 3945 640
rect 3595 615 3945 630
rect -5 600 45 615
rect 95 600 145 615
rect 195 600 245 615
rect 295 600 345 615
rect 395 600 445 615
rect 495 600 545 615
rect 695 600 745 615
rect 795 600 845 615
rect 895 600 945 615
rect 995 600 1045 615
rect 1095 600 1145 615
rect 1195 600 1245 615
rect 1395 600 1445 615
rect 1495 600 1545 615
rect 1595 600 1645 615
rect 1695 600 1745 615
rect 1795 600 1845 615
rect 1895 600 1945 615
rect 2095 600 2145 615
rect 2195 600 2245 615
rect 2295 600 2345 615
rect 2395 600 2445 615
rect 2495 600 2545 615
rect 2595 600 2645 615
rect 2795 600 2845 615
rect 2895 600 2945 615
rect 2995 600 3045 615
rect 3095 600 3145 615
rect 3195 600 3245 615
rect 3295 600 3345 615
rect 3495 600 3545 615
rect 3595 600 3645 615
rect 3695 600 3745 615
rect 3795 600 3845 615
rect 3895 600 3945 615
rect 3995 600 4045 615
rect 4195 600 4245 615
rect 4295 600 4345 640
rect 4395 630 4445 640
rect 4695 640 4995 655
rect 4695 630 4745 640
rect 4395 615 4745 630
rect 4395 600 4445 615
rect 4495 600 4545 615
rect 4595 600 4645 615
rect 4695 600 4745 615
rect 4795 600 4845 640
rect 4895 600 4945 615
rect -5 -15 45 0
rect 95 -15 145 0
rect 195 -15 245 0
rect 295 -15 345 0
rect 395 -15 445 0
rect 495 -15 545 0
rect 695 -15 745 0
rect 795 -15 845 0
rect 895 -15 945 0
rect 995 -15 1045 0
rect 1095 -15 1145 0
rect 1195 -15 1245 0
rect 1395 -15 1445 0
rect 1495 -15 1545 0
rect 1595 -15 1645 0
rect 1695 -15 1745 0
rect 1795 -15 1845 0
rect 1895 -15 1945 0
rect 2095 -15 2145 0
rect 2195 -15 2245 0
rect 2295 -15 2345 0
rect 2395 -15 2445 0
rect 2495 -15 2545 0
rect 2595 -15 2645 0
rect 2795 -15 2845 0
rect 2895 -15 2945 0
rect 2995 -15 3045 0
rect 3095 -15 3145 0
rect 3195 -15 3245 0
rect 3295 -15 3345 0
rect 3495 -15 3545 0
rect 3595 -15 3645 0
rect 3695 -15 3745 0
rect 3795 -15 3845 0
rect 3895 -15 3945 0
rect 3995 -15 4045 0
rect 4195 -15 4245 0
rect 4295 -15 4345 0
rect 4395 -15 4445 0
rect 4495 -15 4545 0
rect 4595 -15 4645 0
rect 4695 -15 4745 0
rect 4795 -15 4845 0
rect -50 -25 45 -15
rect -50 -45 -40 -25
rect -20 -45 45 -25
rect 495 -25 745 -15
rect 495 -30 610 -25
rect -50 -55 45 -45
rect 95 -55 445 -40
rect 600 -45 610 -30
rect 630 -30 745 -25
rect 1195 -25 1445 -15
rect 1195 -30 1310 -25
rect 630 -45 640 -30
rect 600 -55 640 -45
rect 795 -55 1145 -40
rect 1300 -45 1310 -30
rect 1330 -30 1445 -25
rect 1895 -25 2145 -15
rect 1895 -30 2010 -25
rect 1330 -45 1340 -30
rect 1300 -55 1340 -45
rect 1495 -55 1845 -40
rect 2000 -45 2010 -30
rect 2030 -30 2145 -25
rect 2595 -25 2845 -15
rect 2595 -30 2710 -25
rect 2030 -45 2040 -30
rect 2000 -55 2040 -45
rect 2195 -55 2545 -40
rect 2700 -45 2710 -30
rect 2730 -30 2845 -25
rect 3295 -25 3545 -15
rect 3295 -30 3410 -25
rect 2730 -45 2740 -30
rect 2700 -55 2740 -45
rect 2895 -55 3245 -40
rect 3400 -45 3410 -30
rect 3430 -30 3545 -25
rect 3995 -25 4245 -15
rect 3995 -30 4110 -25
rect 3430 -45 3440 -30
rect 3400 -55 3440 -45
rect 3595 -55 3945 -40
rect 4100 -45 4110 -30
rect 4130 -30 4245 -25
rect 4895 -20 4945 0
rect 4895 -30 4990 -20
rect 4130 -45 4140 -30
rect 4100 -55 4140 -45
rect 4295 -55 4645 -40
rect -5 -95 45 -80
rect 95 -95 145 -55
rect 195 -95 245 -80
rect 295 -95 345 -80
rect 395 -95 445 -55
rect 495 -95 545 -80
rect 695 -95 745 -80
rect 795 -95 845 -55
rect 895 -95 945 -80
rect 995 -95 1045 -80
rect 1095 -95 1145 -55
rect 1195 -95 1245 -80
rect 1395 -95 1445 -80
rect 1495 -95 1545 -55
rect 1595 -95 1645 -80
rect 1695 -95 1745 -80
rect 1795 -95 1845 -55
rect 1895 -95 1945 -80
rect 2095 -95 2145 -80
rect 2195 -95 2245 -55
rect 2295 -95 2345 -80
rect 2395 -95 2445 -80
rect 2495 -95 2545 -55
rect 2595 -95 2645 -80
rect 2795 -95 2845 -80
rect 2895 -95 2945 -55
rect 2995 -95 3045 -80
rect 3095 -95 3145 -80
rect 3195 -95 3245 -55
rect 3295 -95 3345 -80
rect 3495 -95 3545 -80
rect 3595 -95 3645 -55
rect 3695 -95 3745 -80
rect 3795 -95 3845 -80
rect 3895 -95 3945 -55
rect 3995 -95 4045 -80
rect 4195 -95 4245 -80
rect 4295 -95 4345 -55
rect 4395 -95 4445 -80
rect 4495 -95 4545 -80
rect 4595 -95 4645 -55
rect 4895 -50 4960 -30
rect 4980 -50 4990 -30
rect 4895 -60 4990 -50
rect 4695 -95 4745 -80
rect -5 -710 45 -695
rect -50 -720 45 -710
rect -50 -740 -40 -720
rect -20 -740 45 -720
rect -50 -750 45 -740
rect 95 -710 145 -695
rect 195 -710 245 -695
rect 295 -710 345 -695
rect 395 -710 445 -695
rect 495 -710 545 -695
rect 695 -710 745 -695
rect 95 -835 110 -710
rect 195 -725 345 -710
rect 495 -720 745 -710
rect 495 -725 610 -720
rect 195 -835 210 -725
rect 600 -740 610 -725
rect 630 -725 745 -720
rect 630 -740 640 -725
rect 690 -730 745 -725
rect 795 -710 845 -695
rect 895 -710 945 -695
rect 995 -710 1045 -695
rect 1095 -710 1145 -695
rect 1195 -710 1245 -695
rect 1395 -710 1445 -695
rect 600 -750 640 -740
rect 795 -835 810 -710
rect 895 -725 1045 -710
rect 1195 -720 1445 -710
rect 1195 -725 1310 -720
rect 895 -835 910 -725
rect 1300 -740 1310 -725
rect 1330 -725 1445 -720
rect 1330 -740 1340 -725
rect 1390 -730 1445 -725
rect 1495 -710 1545 -695
rect 1595 -710 1645 -695
rect 1695 -710 1745 -695
rect 1795 -710 1845 -695
rect 1895 -710 1945 -695
rect 2095 -710 2145 -695
rect 1300 -750 1340 -740
rect 1495 -835 1510 -710
rect 1595 -725 1745 -710
rect 1895 -720 2145 -710
rect 1895 -725 2010 -720
rect 1595 -835 1610 -725
rect 2000 -740 2010 -725
rect 2030 -725 2145 -720
rect 2030 -740 2040 -725
rect 2090 -730 2145 -725
rect 2195 -710 2245 -695
rect 2295 -710 2345 -695
rect 2395 -710 2445 -695
rect 2495 -710 2545 -695
rect 2595 -710 2645 -695
rect 2795 -710 2845 -695
rect 2000 -750 2040 -740
rect 2195 -835 2210 -710
rect 2295 -725 2445 -710
rect 2595 -720 2845 -710
rect 2595 -725 2710 -720
rect 2295 -835 2310 -725
rect 2700 -740 2710 -725
rect 2730 -725 2845 -720
rect 2730 -740 2740 -725
rect 2790 -730 2845 -725
rect 2895 -710 2945 -695
rect 2995 -710 3045 -695
rect 3095 -710 3145 -695
rect 3195 -710 3245 -695
rect 3295 -710 3345 -695
rect 3495 -710 3545 -695
rect 2700 -750 2740 -740
rect 2895 -835 2910 -710
rect 2995 -725 3145 -710
rect 3295 -720 3545 -710
rect 3295 -725 3410 -720
rect 2995 -835 3010 -725
rect 3400 -740 3410 -725
rect 3430 -725 3545 -720
rect 3430 -740 3440 -725
rect 3490 -730 3545 -725
rect 3595 -710 3645 -695
rect 3695 -710 3745 -695
rect 3795 -710 3845 -695
rect 3895 -710 3945 -695
rect 3995 -710 4045 -695
rect 4195 -710 4245 -695
rect 3400 -750 3440 -740
rect 3595 -835 3610 -710
rect 3695 -725 3845 -710
rect 3995 -720 4245 -710
rect 3995 -725 4110 -720
rect 3695 -835 3710 -725
rect 4100 -740 4110 -725
rect 4130 -725 4245 -720
rect 4130 -740 4140 -725
rect 4190 -730 4245 -725
rect 4295 -710 4345 -695
rect 4395 -710 4445 -695
rect 4495 -710 4545 -695
rect 4595 -710 4645 -695
rect 4695 -710 4745 -695
rect 4100 -750 4140 -740
rect 4295 -835 4310 -710
rect 4395 -725 4545 -710
rect 4690 -720 4995 -710
rect 4395 -835 4410 -725
rect 4690 -740 4700 -720
rect 4720 -725 4995 -720
rect 4720 -740 4735 -725
rect 4690 -745 4735 -740
rect 4690 -750 4730 -745
<< polycont >>
rect -40 -45 -20 -25
rect 610 -45 630 -25
rect 1310 -45 1330 -25
rect 2010 -45 2030 -25
rect 2710 -45 2730 -25
rect 3410 -45 3430 -25
rect 4110 -45 4130 -25
rect 4960 -50 4980 -30
rect -40 -740 -20 -720
rect 610 -740 630 -720
rect 1310 -740 1330 -720
rect 2010 -740 2030 -720
rect 2710 -740 2730 -720
rect 3410 -740 3430 -720
rect 4110 -740 4130 -720
rect 4700 -740 4720 -720
<< locali >>
rect 70 685 490 695
rect 70 675 460 685
rect -50 595 -10 600
rect 70 595 90 675
rect 450 665 460 675
rect 480 665 490 685
rect 450 655 490 665
rect 770 685 1190 695
rect 770 675 1160 685
rect 150 645 190 655
rect 150 625 160 645
rect 180 635 190 645
rect 180 625 370 635
rect 150 615 370 625
rect 170 595 190 615
rect 350 595 370 615
rect 450 595 470 655
rect 770 595 790 675
rect 1150 665 1160 675
rect 1180 665 1190 685
rect 1150 655 1190 665
rect 1470 685 1890 695
rect 1470 675 1860 685
rect 850 645 890 655
rect 850 625 860 645
rect 880 635 890 645
rect 880 625 1070 635
rect 850 615 1070 625
rect 870 595 890 615
rect 1050 595 1070 615
rect 1150 595 1170 655
rect 1470 595 1490 675
rect 1850 665 1860 675
rect 1880 665 1890 685
rect 1850 655 1890 665
rect 2170 685 2590 695
rect 2170 675 2560 685
rect 1550 645 1590 655
rect 1550 625 1560 645
rect 1580 635 1590 645
rect 1580 625 1770 635
rect 1550 615 1770 625
rect 1570 595 1590 615
rect 1750 595 1770 615
rect 1850 595 1870 655
rect 2170 595 2190 675
rect 2550 665 2560 675
rect 2580 665 2590 685
rect 2550 655 2590 665
rect 2870 685 3290 695
rect 2870 675 3260 685
rect 2250 645 2290 655
rect 2250 625 2260 645
rect 2280 635 2290 645
rect 2280 625 2470 635
rect 2250 615 2470 625
rect 2270 595 2290 615
rect 2450 595 2470 615
rect 2550 595 2570 655
rect 2870 595 2890 675
rect 3250 665 3260 675
rect 3280 665 3290 685
rect 3250 655 3290 665
rect 3570 685 3990 695
rect 3570 675 3960 685
rect 2950 645 2990 655
rect 2950 625 2960 645
rect 2980 635 2990 645
rect 2980 625 3170 635
rect 2950 615 3170 625
rect 2970 595 2990 615
rect 3150 595 3170 615
rect 3250 595 3270 655
rect 3570 595 3590 675
rect 3950 665 3960 675
rect 3980 665 3990 685
rect 3950 655 3990 665
rect 4370 685 4790 695
rect 4370 675 4760 685
rect 3650 645 3690 655
rect 3650 625 3660 645
rect 3680 635 3690 645
rect 3680 625 3870 635
rect 3650 615 3870 625
rect 3670 595 3690 615
rect 3850 595 3870 615
rect 3950 595 3970 655
rect 4370 595 4390 675
rect 4750 665 4760 675
rect 4780 665 4790 685
rect 4750 655 4790 665
rect 4450 645 4490 655
rect 4450 625 4460 645
rect 4480 635 4490 645
rect 4480 625 4670 635
rect 4450 615 4670 625
rect 4470 595 4490 615
rect 4650 595 4670 615
rect 4750 595 4770 655
rect -100 585 -10 595
rect -100 310 -90 585
rect -70 310 -40 585
rect -20 310 -10 585
rect -100 290 -10 310
rect -100 15 -90 290
rect -70 15 -40 290
rect -20 15 -10 290
rect -100 5 -10 15
rect 50 585 90 595
rect 50 310 60 585
rect 80 310 90 585
rect 50 290 90 310
rect 50 15 60 290
rect 80 15 90 290
rect 50 5 90 15
rect 150 585 190 595
rect 150 310 160 585
rect 180 310 190 585
rect 150 290 190 310
rect 150 15 160 290
rect 180 15 190 290
rect 150 5 190 15
rect 250 585 290 595
rect 250 310 260 585
rect 280 310 290 585
rect 250 290 290 310
rect 250 15 260 290
rect 280 15 290 290
rect 250 5 290 15
rect 350 585 390 595
rect 350 310 360 585
rect 380 310 390 585
rect 350 290 390 310
rect 350 15 360 290
rect 380 15 390 290
rect 350 5 390 15
rect 450 585 490 595
rect 450 310 460 585
rect 480 310 490 585
rect 450 290 490 310
rect 450 15 460 290
rect 480 15 490 290
rect 450 5 490 15
rect 550 585 690 595
rect 550 310 560 585
rect 580 310 610 585
rect 630 310 660 585
rect 680 310 690 585
rect 550 290 690 310
rect 550 15 560 290
rect 580 15 610 290
rect 630 15 660 290
rect 680 15 690 290
rect 550 5 690 15
rect 750 585 790 595
rect 750 310 760 585
rect 780 310 790 585
rect 750 290 790 310
rect 750 15 760 290
rect 780 15 790 290
rect 750 5 790 15
rect 850 585 890 595
rect 850 310 860 585
rect 880 310 890 585
rect 850 290 890 310
rect 850 15 860 290
rect 880 15 890 290
rect 850 5 890 15
rect 950 585 990 595
rect 950 310 960 585
rect 980 310 990 585
rect 950 290 990 310
rect 950 15 960 290
rect 980 15 990 290
rect 950 5 990 15
rect 1050 585 1090 595
rect 1050 310 1060 585
rect 1080 310 1090 585
rect 1050 290 1090 310
rect 1050 15 1060 290
rect 1080 15 1090 290
rect 1050 5 1090 15
rect 1150 585 1190 595
rect 1150 310 1160 585
rect 1180 310 1190 585
rect 1150 290 1190 310
rect 1150 15 1160 290
rect 1180 15 1190 290
rect 1150 5 1190 15
rect 1250 585 1390 595
rect 1250 310 1260 585
rect 1280 310 1310 585
rect 1330 310 1360 585
rect 1380 310 1390 585
rect 1250 290 1390 310
rect 1250 15 1260 290
rect 1280 15 1310 290
rect 1330 15 1360 290
rect 1380 15 1390 290
rect 1250 5 1390 15
rect 1450 585 1490 595
rect 1450 310 1460 585
rect 1480 310 1490 585
rect 1450 290 1490 310
rect 1450 15 1460 290
rect 1480 15 1490 290
rect 1450 5 1490 15
rect 1550 585 1590 595
rect 1550 310 1560 585
rect 1580 310 1590 585
rect 1550 290 1590 310
rect 1550 15 1560 290
rect 1580 15 1590 290
rect 1550 5 1590 15
rect 1650 585 1690 595
rect 1650 310 1660 585
rect 1680 310 1690 585
rect 1650 290 1690 310
rect 1650 15 1660 290
rect 1680 15 1690 290
rect 1650 5 1690 15
rect 1750 585 1790 595
rect 1750 310 1760 585
rect 1780 310 1790 585
rect 1750 290 1790 310
rect 1750 15 1760 290
rect 1780 15 1790 290
rect 1750 5 1790 15
rect 1850 585 1890 595
rect 1850 310 1860 585
rect 1880 310 1890 585
rect 1850 290 1890 310
rect 1850 15 1860 290
rect 1880 15 1890 290
rect 1850 5 1890 15
rect 1950 585 2090 595
rect 1950 310 1960 585
rect 1980 310 2010 585
rect 2030 310 2060 585
rect 2080 310 2090 585
rect 1950 290 2090 310
rect 1950 15 1960 290
rect 1980 15 2010 290
rect 2030 15 2060 290
rect 2080 15 2090 290
rect 1950 5 2090 15
rect 2150 585 2190 595
rect 2150 310 2160 585
rect 2180 310 2190 585
rect 2150 290 2190 310
rect 2150 15 2160 290
rect 2180 15 2190 290
rect 2150 5 2190 15
rect 2250 585 2290 595
rect 2250 310 2260 585
rect 2280 310 2290 585
rect 2250 290 2290 310
rect 2250 15 2260 290
rect 2280 15 2290 290
rect 2250 5 2290 15
rect 2350 585 2390 595
rect 2350 310 2360 585
rect 2380 310 2390 585
rect 2350 290 2390 310
rect 2350 15 2360 290
rect 2380 15 2390 290
rect 2350 5 2390 15
rect 2450 585 2490 595
rect 2450 310 2460 585
rect 2480 310 2490 585
rect 2450 290 2490 310
rect 2450 15 2460 290
rect 2480 15 2490 290
rect 2450 5 2490 15
rect 2550 585 2590 595
rect 2550 310 2560 585
rect 2580 310 2590 585
rect 2550 290 2590 310
rect 2550 15 2560 290
rect 2580 15 2590 290
rect 2550 5 2590 15
rect 2650 585 2790 595
rect 2650 310 2660 585
rect 2680 310 2710 585
rect 2730 310 2760 585
rect 2780 310 2790 585
rect 2650 290 2790 310
rect 2650 15 2660 290
rect 2680 15 2710 290
rect 2730 15 2760 290
rect 2780 15 2790 290
rect 2650 5 2790 15
rect 2850 585 2890 595
rect 2850 310 2860 585
rect 2880 310 2890 585
rect 2850 290 2890 310
rect 2850 15 2860 290
rect 2880 15 2890 290
rect 2850 5 2890 15
rect 2950 585 2990 595
rect 2950 310 2960 585
rect 2980 310 2990 585
rect 2950 290 2990 310
rect 2950 15 2960 290
rect 2980 15 2990 290
rect 2950 5 2990 15
rect 3050 585 3090 595
rect 3050 310 3060 585
rect 3080 310 3090 585
rect 3050 290 3090 310
rect 3050 15 3060 290
rect 3080 15 3090 290
rect 3050 5 3090 15
rect 3150 585 3190 595
rect 3150 310 3160 585
rect 3180 310 3190 585
rect 3150 290 3190 310
rect 3150 15 3160 290
rect 3180 15 3190 290
rect 3150 5 3190 15
rect 3250 585 3290 595
rect 3250 310 3260 585
rect 3280 310 3290 585
rect 3250 290 3290 310
rect 3250 15 3260 290
rect 3280 15 3290 290
rect 3250 5 3290 15
rect 3350 585 3490 595
rect 3350 310 3360 585
rect 3380 310 3410 585
rect 3430 310 3460 585
rect 3480 310 3490 585
rect 3350 290 3490 310
rect 3350 15 3360 290
rect 3380 15 3410 290
rect 3430 15 3460 290
rect 3480 15 3490 290
rect 3350 5 3490 15
rect 3550 585 3590 595
rect 3550 310 3560 585
rect 3580 310 3590 585
rect 3550 290 3590 310
rect 3550 15 3560 290
rect 3580 15 3590 290
rect 3550 5 3590 15
rect 3650 585 3690 595
rect 3650 310 3660 585
rect 3680 310 3690 585
rect 3650 290 3690 310
rect 3650 15 3660 290
rect 3680 15 3690 290
rect 3650 5 3690 15
rect 3750 585 3790 595
rect 3750 310 3760 585
rect 3780 310 3790 585
rect 3750 290 3790 310
rect 3750 15 3760 290
rect 3780 15 3790 290
rect 3750 5 3790 15
rect 3850 585 3890 595
rect 3850 310 3860 585
rect 3880 310 3890 585
rect 3850 290 3890 310
rect 3850 15 3860 290
rect 3880 15 3890 290
rect 3850 5 3890 15
rect 3950 585 3990 595
rect 3950 310 3960 585
rect 3980 310 3990 585
rect 3950 290 3990 310
rect 3950 15 3960 290
rect 3980 15 3990 290
rect 3950 5 3990 15
rect 4050 585 4190 595
rect 4050 310 4060 585
rect 4080 310 4110 585
rect 4130 310 4160 585
rect 4180 310 4190 585
rect 4050 290 4190 310
rect 4050 15 4060 290
rect 4080 15 4110 290
rect 4130 15 4160 290
rect 4180 15 4190 290
rect 4050 5 4190 15
rect 4250 585 4290 595
rect 4250 310 4260 585
rect 4280 310 4290 585
rect 4250 290 4290 310
rect 4250 15 4260 290
rect 4280 15 4290 290
rect 4250 5 4290 15
rect 4350 585 4390 595
rect 4350 310 4360 585
rect 4380 310 4390 585
rect 4350 290 4390 310
rect 4350 15 4360 290
rect 4380 15 4390 290
rect 4350 5 4390 15
rect 4450 585 4490 595
rect 4450 310 4460 585
rect 4480 310 4490 585
rect 4450 290 4490 310
rect 4450 15 4460 290
rect 4480 15 4490 290
rect 4450 5 4490 15
rect 4550 585 4590 595
rect 4550 310 4560 585
rect 4580 310 4590 585
rect 4550 290 4590 310
rect 4550 15 4560 290
rect 4580 15 4590 290
rect 4550 5 4590 15
rect 4650 585 4690 595
rect 4650 310 4660 585
rect 4680 310 4690 585
rect 4650 290 4690 310
rect 4650 15 4660 290
rect 4680 15 4690 290
rect 4650 5 4690 15
rect 4750 585 4790 595
rect 4750 310 4760 585
rect 4780 310 4790 585
rect 4750 290 4790 310
rect 4750 15 4760 290
rect 4780 15 4790 290
rect 4750 5 4790 15
rect 4850 585 4890 595
rect 4850 310 4860 585
rect 4880 310 4890 585
rect 4850 290 4890 310
rect 4850 15 4860 290
rect 4880 15 4890 290
rect 4850 5 4890 15
rect 4950 585 4990 595
rect 4950 310 4960 585
rect 4980 310 4990 585
rect 4950 290 4990 310
rect 4950 15 4960 290
rect 4980 15 4990 290
rect -50 -25 -10 5
rect -50 -45 -40 -25
rect -20 -45 -10 -25
rect -50 -55 -10 -45
rect 260 -60 280 5
rect 550 0 590 5
rect 570 -15 590 0
rect 650 0 690 5
rect 650 -15 670 0
rect 570 -25 670 -15
rect 570 -35 610 -25
rect 600 -45 610 -35
rect 630 -35 670 -25
rect 630 -45 640 -35
rect 600 -55 640 -45
rect 960 -60 980 5
rect 1250 0 1290 5
rect 1270 -15 1290 0
rect 1350 0 1390 5
rect 1350 -15 1370 0
rect 1270 -25 1370 -15
rect 1270 -35 1310 -25
rect 1300 -45 1310 -35
rect 1330 -35 1370 -25
rect 1330 -45 1340 -35
rect 1300 -55 1340 -45
rect 1660 -60 1680 5
rect 1950 0 1990 5
rect 1970 -15 1990 0
rect 2050 0 2090 5
rect 2050 -15 2070 0
rect 1970 -25 2070 -15
rect 1970 -35 2010 -25
rect 2000 -45 2010 -35
rect 2030 -35 2070 -25
rect 2030 -45 2040 -35
rect 2000 -55 2040 -45
rect 2360 -60 2380 5
rect 2650 0 2690 5
rect 2670 -15 2690 0
rect 2750 0 2790 5
rect 2750 -15 2770 0
rect 2670 -25 2770 -15
rect 2670 -35 2710 -25
rect 2700 -45 2710 -35
rect 2730 -35 2770 -25
rect 2730 -45 2740 -35
rect 2700 -55 2740 -45
rect 3060 -60 3080 5
rect 3350 0 3390 5
rect 3370 -15 3390 0
rect 3450 0 3490 5
rect 3450 -15 3470 0
rect 3370 -25 3470 -15
rect 3370 -35 3410 -25
rect 3400 -45 3410 -35
rect 3430 -35 3470 -25
rect 3430 -45 3440 -35
rect 3400 -55 3440 -45
rect 3760 -60 3780 5
rect 4050 0 4090 5
rect 4070 -15 4090 0
rect 4150 0 4190 5
rect 4150 -15 4170 0
rect 4070 -25 4170 -15
rect 4560 -20 4580 5
rect 4950 0 4990 15
rect 4970 -20 4990 0
rect 4070 -35 4110 -25
rect 4100 -45 4110 -35
rect 4130 -35 4170 -25
rect 4130 -45 4140 -35
rect 4100 -55 4140 -45
rect 4460 -40 4580 -20
rect 4950 -30 4990 -20
rect 4460 -60 4480 -40
rect 4950 -50 4960 -30
rect 4980 -50 4990 -30
rect 4950 -60 4990 -50
rect 170 -80 370 -60
rect 170 -100 190 -80
rect 350 -100 370 -80
rect 870 -80 1070 -60
rect 870 -100 890 -80
rect 1050 -100 1070 -80
rect 1570 -80 1770 -60
rect 1570 -100 1590 -80
rect 1750 -100 1770 -80
rect 2270 -80 2470 -60
rect 2270 -100 2290 -80
rect 2450 -100 2470 -80
rect 2970 -80 3170 -60
rect 2970 -100 2990 -80
rect 3150 -100 3170 -80
rect 3670 -80 3870 -60
rect 3670 -100 3690 -80
rect 3850 -100 3870 -80
rect 4370 -80 4570 -60
rect 4370 -100 4390 -80
rect 4550 -100 4570 -80
rect -100 -110 -10 -100
rect -100 -385 -90 -110
rect -70 -385 -40 -110
rect -20 -385 -10 -110
rect -100 -405 -10 -385
rect -100 -680 -90 -405
rect -70 -680 -40 -405
rect -20 -680 -10 -405
rect -100 -690 -10 -680
rect 50 -110 90 -100
rect 50 -385 60 -110
rect 80 -385 90 -110
rect 50 -405 90 -385
rect 50 -680 60 -405
rect 80 -680 90 -405
rect 50 -690 90 -680
rect 150 -110 190 -100
rect 150 -385 160 -110
rect 180 -385 190 -110
rect 150 -405 190 -385
rect 150 -680 160 -405
rect 180 -680 190 -405
rect 150 -690 190 -680
rect 250 -110 290 -100
rect 250 -385 260 -110
rect 280 -385 290 -110
rect 250 -405 290 -385
rect 250 -680 260 -405
rect 280 -680 290 -405
rect 250 -690 290 -680
rect 350 -110 390 -100
rect 350 -385 360 -110
rect 380 -385 390 -110
rect 350 -405 390 -385
rect 350 -680 360 -405
rect 380 -680 390 -405
rect 350 -690 390 -680
rect 450 -110 490 -100
rect 450 -385 460 -110
rect 480 -385 490 -110
rect 450 -405 490 -385
rect 450 -680 460 -405
rect 480 -680 490 -405
rect 450 -690 490 -680
rect 550 -110 690 -100
rect 550 -385 560 -110
rect 580 -385 610 -110
rect 630 -385 660 -110
rect 680 -385 690 -110
rect 550 -405 690 -385
rect 550 -680 560 -405
rect 580 -680 610 -405
rect 630 -680 660 -405
rect 680 -680 690 -405
rect 550 -690 690 -680
rect 750 -110 790 -100
rect 750 -385 760 -110
rect 780 -385 790 -110
rect 750 -405 790 -385
rect 750 -680 760 -405
rect 780 -680 790 -405
rect 750 -690 790 -680
rect 850 -110 890 -100
rect 850 -385 860 -110
rect 880 -385 890 -110
rect 850 -405 890 -385
rect 850 -680 860 -405
rect 880 -680 890 -405
rect 850 -690 890 -680
rect 950 -110 990 -100
rect 950 -385 960 -110
rect 980 -385 990 -110
rect 950 -405 990 -385
rect 950 -680 960 -405
rect 980 -680 990 -405
rect 950 -690 990 -680
rect 1050 -110 1090 -100
rect 1050 -385 1060 -110
rect 1080 -385 1090 -110
rect 1050 -405 1090 -385
rect 1050 -680 1060 -405
rect 1080 -680 1090 -405
rect 1050 -690 1090 -680
rect 1150 -110 1190 -100
rect 1150 -385 1160 -110
rect 1180 -385 1190 -110
rect 1150 -405 1190 -385
rect 1150 -680 1160 -405
rect 1180 -680 1190 -405
rect 1150 -690 1190 -680
rect 1250 -110 1390 -100
rect 1250 -385 1260 -110
rect 1280 -385 1310 -110
rect 1330 -385 1360 -110
rect 1380 -385 1390 -110
rect 1250 -405 1390 -385
rect 1250 -680 1260 -405
rect 1280 -680 1310 -405
rect 1330 -680 1360 -405
rect 1380 -680 1390 -405
rect 1250 -690 1390 -680
rect 1450 -110 1490 -100
rect 1450 -385 1460 -110
rect 1480 -385 1490 -110
rect 1450 -405 1490 -385
rect 1450 -680 1460 -405
rect 1480 -680 1490 -405
rect 1450 -690 1490 -680
rect 1550 -110 1590 -100
rect 1550 -385 1560 -110
rect 1580 -385 1590 -110
rect 1550 -405 1590 -385
rect 1550 -680 1560 -405
rect 1580 -680 1590 -405
rect 1550 -690 1590 -680
rect 1650 -110 1690 -100
rect 1650 -385 1660 -110
rect 1680 -385 1690 -110
rect 1650 -405 1690 -385
rect 1650 -680 1660 -405
rect 1680 -680 1690 -405
rect 1650 -690 1690 -680
rect 1750 -110 1790 -100
rect 1750 -385 1760 -110
rect 1780 -385 1790 -110
rect 1750 -405 1790 -385
rect 1750 -680 1760 -405
rect 1780 -680 1790 -405
rect 1750 -690 1790 -680
rect 1850 -110 1890 -100
rect 1850 -385 1860 -110
rect 1880 -385 1890 -110
rect 1850 -405 1890 -385
rect 1850 -680 1860 -405
rect 1880 -680 1890 -405
rect 1850 -690 1890 -680
rect 1950 -110 2090 -100
rect 1950 -385 1960 -110
rect 1980 -385 2010 -110
rect 2030 -385 2060 -110
rect 2080 -385 2090 -110
rect 1950 -405 2090 -385
rect 1950 -680 1960 -405
rect 1980 -680 2010 -405
rect 2030 -680 2060 -405
rect 2080 -680 2090 -405
rect 1950 -690 2090 -680
rect 2150 -110 2190 -100
rect 2150 -385 2160 -110
rect 2180 -385 2190 -110
rect 2150 -405 2190 -385
rect 2150 -680 2160 -405
rect 2180 -680 2190 -405
rect 2150 -690 2190 -680
rect 2250 -110 2290 -100
rect 2250 -385 2260 -110
rect 2280 -385 2290 -110
rect 2250 -405 2290 -385
rect 2250 -680 2260 -405
rect 2280 -680 2290 -405
rect 2250 -690 2290 -680
rect 2350 -110 2390 -100
rect 2350 -385 2360 -110
rect 2380 -385 2390 -110
rect 2350 -405 2390 -385
rect 2350 -680 2360 -405
rect 2380 -680 2390 -405
rect 2350 -690 2390 -680
rect 2450 -110 2490 -100
rect 2450 -385 2460 -110
rect 2480 -385 2490 -110
rect 2450 -405 2490 -385
rect 2450 -680 2460 -405
rect 2480 -680 2490 -405
rect 2450 -690 2490 -680
rect 2550 -110 2590 -100
rect 2550 -385 2560 -110
rect 2580 -385 2590 -110
rect 2550 -405 2590 -385
rect 2550 -680 2560 -405
rect 2580 -680 2590 -405
rect 2550 -690 2590 -680
rect 2650 -110 2790 -100
rect 2650 -385 2660 -110
rect 2680 -385 2710 -110
rect 2730 -385 2760 -110
rect 2780 -385 2790 -110
rect 2650 -405 2790 -385
rect 2650 -680 2660 -405
rect 2680 -680 2710 -405
rect 2730 -680 2760 -405
rect 2780 -680 2790 -405
rect 2650 -690 2790 -680
rect 2850 -110 2890 -100
rect 2850 -385 2860 -110
rect 2880 -385 2890 -110
rect 2850 -405 2890 -385
rect 2850 -680 2860 -405
rect 2880 -680 2890 -405
rect 2850 -690 2890 -680
rect 2950 -110 2990 -100
rect 2950 -385 2960 -110
rect 2980 -385 2990 -110
rect 2950 -405 2990 -385
rect 2950 -680 2960 -405
rect 2980 -680 2990 -405
rect 2950 -690 2990 -680
rect 3050 -110 3090 -100
rect 3050 -385 3060 -110
rect 3080 -385 3090 -110
rect 3050 -405 3090 -385
rect 3050 -680 3060 -405
rect 3080 -680 3090 -405
rect 3050 -690 3090 -680
rect 3150 -110 3190 -100
rect 3150 -385 3160 -110
rect 3180 -385 3190 -110
rect 3150 -405 3190 -385
rect 3150 -680 3160 -405
rect 3180 -680 3190 -405
rect 3150 -690 3190 -680
rect 3250 -110 3290 -100
rect 3250 -385 3260 -110
rect 3280 -385 3290 -110
rect 3250 -405 3290 -385
rect 3250 -680 3260 -405
rect 3280 -680 3290 -405
rect 3250 -690 3290 -680
rect 3350 -110 3490 -100
rect 3350 -385 3360 -110
rect 3380 -385 3410 -110
rect 3430 -385 3460 -110
rect 3480 -385 3490 -110
rect 3350 -405 3490 -385
rect 3350 -680 3360 -405
rect 3380 -680 3410 -405
rect 3430 -680 3460 -405
rect 3480 -680 3490 -405
rect 3350 -690 3490 -680
rect 3550 -110 3590 -100
rect 3550 -385 3560 -110
rect 3580 -385 3590 -110
rect 3550 -405 3590 -385
rect 3550 -680 3560 -405
rect 3580 -680 3590 -405
rect 3550 -690 3590 -680
rect 3650 -110 3690 -100
rect 3650 -385 3660 -110
rect 3680 -385 3690 -110
rect 3650 -405 3690 -385
rect 3650 -680 3660 -405
rect 3680 -680 3690 -405
rect 3650 -690 3690 -680
rect 3750 -110 3790 -100
rect 3750 -385 3760 -110
rect 3780 -385 3790 -110
rect 3750 -405 3790 -385
rect 3750 -680 3760 -405
rect 3780 -680 3790 -405
rect 3750 -690 3790 -680
rect 3850 -110 3890 -100
rect 3850 -385 3860 -110
rect 3880 -385 3890 -110
rect 3850 -405 3890 -385
rect 3850 -680 3860 -405
rect 3880 -680 3890 -405
rect 3850 -690 3890 -680
rect 3950 -110 3990 -100
rect 3950 -385 3960 -110
rect 3980 -385 3990 -110
rect 3950 -405 3990 -385
rect 3950 -680 3960 -405
rect 3980 -680 3990 -405
rect 3950 -690 3990 -680
rect 4050 -110 4190 -100
rect 4050 -385 4060 -110
rect 4080 -385 4110 -110
rect 4130 -385 4160 -110
rect 4180 -385 4190 -110
rect 4050 -405 4190 -385
rect 4050 -680 4060 -405
rect 4080 -680 4110 -405
rect 4130 -680 4160 -405
rect 4180 -680 4190 -405
rect 4050 -690 4190 -680
rect 4250 -110 4290 -100
rect 4250 -385 4260 -110
rect 4280 -385 4290 -110
rect 4250 -405 4290 -385
rect 4250 -680 4260 -405
rect 4280 -680 4290 -405
rect 4250 -690 4290 -680
rect 4350 -110 4390 -100
rect 4350 -385 4360 -110
rect 4380 -385 4390 -110
rect 4350 -405 4390 -385
rect 4350 -680 4360 -405
rect 4380 -680 4390 -405
rect 4350 -690 4390 -680
rect 4450 -110 4490 -100
rect 4450 -385 4460 -110
rect 4480 -385 4490 -110
rect 4450 -405 4490 -385
rect 4450 -680 4460 -405
rect 4480 -680 4490 -405
rect 4450 -690 4490 -680
rect 4550 -110 4590 -100
rect 4550 -385 4560 -110
rect 4580 -385 4590 -110
rect 4550 -405 4590 -385
rect 4550 -680 4560 -405
rect 4580 -680 4590 -405
rect 4550 -690 4590 -680
rect 4650 -110 4690 -100
rect 4650 -385 4660 -110
rect 4680 -385 4690 -110
rect 4650 -405 4690 -385
rect 4650 -680 4660 -405
rect 4680 -680 4690 -405
rect 4650 -690 4690 -680
rect 4750 -110 4795 -100
rect 4750 -385 4760 -110
rect 4780 -385 4795 -110
rect 4750 -405 4795 -385
rect 4750 -680 4760 -405
rect 4780 -680 4795 -405
rect 4750 -690 4795 -680
rect -50 -720 -10 -690
rect -50 -740 -40 -720
rect -20 -740 -10 -720
rect -50 -750 -10 -740
rect 70 -770 90 -690
rect 450 -770 470 -690
rect 550 -710 590 -690
rect 650 -710 690 -690
rect 550 -720 690 -710
rect 550 -730 610 -720
rect 600 -740 610 -730
rect 630 -730 690 -720
rect 630 -740 640 -730
rect 600 -750 640 -740
rect 770 -770 790 -690
rect 1150 -770 1170 -690
rect 1250 -710 1290 -690
rect 1350 -710 1390 -690
rect 1250 -720 1390 -710
rect 1250 -730 1310 -720
rect 1300 -740 1310 -730
rect 1330 -730 1390 -720
rect 1330 -740 1340 -730
rect 1300 -750 1340 -740
rect 1470 -770 1490 -690
rect 1850 -770 1870 -690
rect 1950 -710 1990 -690
rect 2050 -710 2090 -690
rect 1950 -720 2090 -710
rect 1950 -730 2010 -720
rect 2000 -740 2010 -730
rect 2030 -730 2090 -720
rect 2030 -740 2040 -730
rect 2000 -750 2040 -740
rect 2170 -770 2190 -690
rect 2550 -770 2570 -690
rect 2650 -710 2690 -690
rect 2750 -710 2790 -690
rect 2650 -720 2790 -710
rect 2650 -730 2710 -720
rect 2700 -740 2710 -730
rect 2730 -730 2790 -720
rect 2730 -740 2740 -730
rect 2700 -750 2740 -740
rect 2870 -770 2890 -690
rect 3250 -770 3270 -690
rect 3350 -710 3390 -690
rect 3450 -710 3490 -690
rect 3350 -720 3490 -710
rect 3350 -730 3410 -720
rect 3400 -740 3410 -730
rect 3430 -730 3490 -720
rect 3430 -740 3440 -730
rect 3400 -750 3440 -740
rect 3570 -770 3590 -690
rect 3950 -770 3970 -690
rect 4050 -710 4090 -690
rect 4150 -710 4190 -690
rect 4050 -720 4190 -710
rect 4050 -730 4110 -720
rect 4100 -740 4110 -730
rect 4130 -730 4190 -720
rect 4130 -740 4140 -730
rect 4100 -750 4140 -740
rect 4270 -770 4290 -690
rect 4650 -770 4670 -690
rect 4750 -710 4790 -690
rect 4690 -720 4995 -710
rect 4690 -740 4700 -720
rect 4720 -730 4995 -720
rect 4720 -740 4730 -730
rect 4690 -750 4730 -740
rect -165 -790 4995 -770
<< viali >>
rect 460 665 480 685
rect 160 625 180 645
rect 1160 665 1180 685
rect 860 625 880 645
rect 1860 665 1880 685
rect 1560 625 1580 645
rect 2560 665 2580 685
rect 2260 625 2280 645
rect 3260 665 3280 685
rect 2960 625 2980 645
rect 3960 665 3980 685
rect 3660 625 3680 645
rect 4760 665 4780 685
rect 4460 625 4480 645
rect -90 310 -70 585
rect -40 310 -20 585
rect -90 15 -70 290
rect -40 15 -20 290
rect 560 310 580 585
rect 610 310 630 585
rect 660 310 680 585
rect 560 15 580 290
rect 610 15 630 290
rect 660 15 680 290
rect 1260 310 1280 585
rect 1310 310 1330 585
rect 1360 310 1380 585
rect 1260 15 1280 290
rect 1310 15 1330 290
rect 1360 15 1380 290
rect 1960 310 1980 585
rect 2010 310 2030 585
rect 2060 310 2080 585
rect 1960 15 1980 290
rect 2010 15 2030 290
rect 2060 15 2080 290
rect 2660 310 2680 585
rect 2710 310 2730 585
rect 2760 310 2780 585
rect 2660 15 2680 290
rect 2710 15 2730 290
rect 2760 15 2780 290
rect 3360 310 3380 585
rect 3410 310 3430 585
rect 3460 310 3480 585
rect 3360 15 3380 290
rect 3410 15 3430 290
rect 3460 15 3480 290
rect 4060 310 4080 585
rect 4110 310 4130 585
rect 4160 310 4180 585
rect 4060 15 4080 290
rect 4110 15 4130 290
rect 4160 15 4180 290
rect 4260 310 4280 585
rect 4260 15 4280 290
rect 4860 310 4880 585
rect 4860 15 4880 290
rect 4960 310 4980 585
rect 4960 15 4980 290
rect -40 -45 -20 -25
rect 610 -45 630 -25
rect 1310 -45 1330 -25
rect 2010 -45 2030 -25
rect 2710 -45 2730 -25
rect 3410 -45 3430 -25
rect 4110 -45 4130 -25
rect 4960 -50 4980 -30
rect -90 -385 -70 -110
rect -40 -385 -20 -110
rect -90 -680 -70 -405
rect -40 -680 -20 -405
rect 260 -385 280 -110
rect 260 -680 280 -405
rect 560 -385 580 -110
rect 610 -385 630 -110
rect 660 -385 680 -110
rect 560 -680 580 -405
rect 610 -680 630 -405
rect 660 -680 680 -405
rect 960 -385 980 -110
rect 960 -680 980 -405
rect 1260 -385 1280 -110
rect 1310 -385 1330 -110
rect 1360 -385 1380 -110
rect 1260 -680 1280 -405
rect 1310 -680 1330 -405
rect 1360 -680 1380 -405
rect 1660 -385 1680 -110
rect 1660 -680 1680 -405
rect 1960 -385 1980 -110
rect 2010 -385 2030 -110
rect 2060 -385 2080 -110
rect 1960 -680 1980 -405
rect 2010 -680 2030 -405
rect 2060 -680 2080 -405
rect 2360 -385 2380 -110
rect 2360 -680 2380 -405
rect 2660 -385 2680 -110
rect 2710 -385 2730 -110
rect 2760 -385 2780 -110
rect 2660 -680 2680 -405
rect 2710 -680 2730 -405
rect 2760 -680 2780 -405
rect 3060 -385 3080 -110
rect 3060 -680 3080 -405
rect 3360 -385 3380 -110
rect 3410 -385 3430 -110
rect 3460 -385 3480 -110
rect 3360 -680 3380 -405
rect 3410 -680 3430 -405
rect 3460 -680 3480 -405
rect 3760 -385 3780 -110
rect 3760 -680 3780 -405
rect 4060 -385 4080 -110
rect 4110 -385 4130 -110
rect 4160 -385 4180 -110
rect 4060 -680 4080 -405
rect 4110 -680 4130 -405
rect 4160 -680 4180 -405
rect 4460 -385 4480 -110
rect 4460 -680 4480 -405
rect 4760 -385 4780 -110
rect 4760 -680 4780 -405
<< metal1 >>
rect -165 655 190 695
rect 450 685 890 695
rect 450 665 460 685
rect 480 665 890 685
rect 450 655 890 665
rect 1150 685 1590 695
rect 1150 665 1160 685
rect 1180 665 1590 685
rect 1150 655 1590 665
rect 1850 685 2290 695
rect 1850 665 1860 685
rect 1880 665 2290 685
rect 1850 655 2290 665
rect 2550 685 2990 695
rect 2550 665 2560 685
rect 2580 665 2990 685
rect 2550 655 2990 665
rect 3250 685 3690 695
rect 3250 665 3260 685
rect 3280 665 3690 685
rect 3250 655 3690 665
rect 3950 685 4490 695
rect 3950 665 3960 685
rect 3980 665 4490 685
rect 3950 655 4490 665
rect 4750 685 4995 695
rect 4750 665 4760 685
rect 4780 665 4995 685
rect 4750 655 4995 665
rect 150 645 190 655
rect 150 625 160 645
rect 180 625 190 645
rect 150 615 190 625
rect 850 645 890 655
rect 850 625 860 645
rect 880 625 890 645
rect 850 615 890 625
rect 1550 645 1590 655
rect 1550 625 1560 645
rect 1580 625 1590 645
rect 1550 615 1590 625
rect 2250 645 2290 655
rect 2250 625 2260 645
rect 2280 625 2290 645
rect 2250 615 2290 625
rect 2950 645 2990 655
rect 2950 625 2960 645
rect 2980 625 2990 645
rect 2950 615 2990 625
rect 3650 645 3690 655
rect 3650 625 3660 645
rect 3680 625 3690 645
rect 3650 615 3690 625
rect 4450 645 4490 655
rect 4450 625 4460 645
rect 4480 625 4490 645
rect 4450 615 4490 625
rect -165 585 120 600
rect 220 585 820 600
rect 920 585 1520 600
rect 1620 585 2220 600
rect 2320 585 2920 600
rect 3020 585 3620 600
rect 3720 585 4420 600
rect 4520 585 4995 600
rect -165 310 -90 585
rect -70 310 -40 585
rect -20 310 560 585
rect 580 310 610 585
rect 630 310 660 585
rect 680 310 1260 585
rect 1280 310 1310 585
rect 1330 310 1360 585
rect 1380 310 1960 585
rect 1980 310 2010 585
rect 2030 310 2060 585
rect 2080 310 2660 585
rect 2680 310 2710 585
rect 2730 310 2760 585
rect 2780 310 3360 585
rect 3380 310 3410 585
rect 3430 310 3460 585
rect 3480 310 4060 585
rect 4080 310 4110 585
rect 4130 310 4160 585
rect 4180 310 4260 585
rect 4280 310 4860 585
rect 4880 310 4960 585
rect 4980 310 4995 585
rect -165 290 4995 310
rect -165 15 -90 290
rect -70 15 -40 290
rect -20 15 560 290
rect 580 15 610 290
rect 630 15 660 290
rect 680 15 1260 290
rect 1280 15 1310 290
rect 1330 15 1360 290
rect 1380 15 1960 290
rect 1980 15 2010 290
rect 2030 15 2060 290
rect 2080 15 2660 290
rect 2680 15 2710 290
rect 2730 15 2760 290
rect 2780 15 3360 290
rect 3380 15 3410 290
rect 3430 15 3460 290
rect 3480 15 4060 290
rect 4080 15 4110 290
rect 4130 15 4160 290
rect 4180 15 4260 290
rect 4280 15 4860 290
rect 4880 15 4960 290
rect 4980 15 4995 290
rect -165 -25 4995 15
rect -165 -45 -40 -25
rect -20 -45 610 -25
rect 630 -45 1310 -25
rect 1330 -45 2010 -25
rect 2030 -45 2710 -25
rect 2730 -45 3410 -25
rect 3430 -45 4110 -25
rect 4130 -30 4995 -25
rect 4130 -45 4960 -30
rect -165 -50 4960 -45
rect 4980 -50 4995 -30
rect -165 -110 4995 -50
rect -165 -385 -90 -110
rect -70 -385 -40 -110
rect -20 -385 260 -110
rect 280 -385 560 -110
rect 580 -385 610 -110
rect 630 -385 660 -110
rect 680 -385 960 -110
rect 980 -385 1260 -110
rect 1280 -385 1310 -110
rect 1330 -385 1360 -110
rect 1380 -385 1660 -110
rect 1680 -385 1960 -110
rect 1980 -385 2010 -110
rect 2030 -385 2060 -110
rect 2080 -385 2360 -110
rect 2380 -385 2660 -110
rect 2680 -385 2710 -110
rect 2730 -385 2760 -110
rect 2780 -385 3060 -110
rect 3080 -385 3360 -110
rect 3380 -385 3410 -110
rect 3430 -385 3460 -110
rect 3480 -385 3760 -110
rect 3780 -385 4060 -110
rect 4080 -385 4110 -110
rect 4130 -385 4160 -110
rect 4180 -385 4460 -110
rect 4480 -385 4760 -110
rect 4780 -385 4995 -110
rect -165 -405 4995 -385
rect -165 -680 -90 -405
rect -70 -680 -40 -405
rect -20 -680 260 -405
rect 280 -680 560 -405
rect 580 -680 610 -405
rect 630 -680 660 -405
rect 680 -680 960 -405
rect 980 -680 1260 -405
rect 1280 -680 1310 -405
rect 1330 -680 1360 -405
rect 1380 -680 1660 -405
rect 1680 -680 1960 -405
rect 1980 -680 2010 -405
rect 2030 -680 2060 -405
rect 2080 -680 2360 -405
rect 2380 -680 2660 -405
rect 2680 -680 2710 -405
rect 2730 -680 2760 -405
rect 2780 -680 3060 -405
rect 3080 -680 3360 -405
rect 3380 -680 3410 -405
rect 3430 -680 3460 -405
rect 3480 -680 3760 -405
rect 3780 -680 4060 -405
rect 4080 -680 4110 -405
rect 4130 -680 4160 -405
rect 4180 -680 4460 -405
rect 4480 -680 4760 -405
rect 4780 -680 4995 -405
rect -165 -695 4995 -680
<< labels >>
rlabel metal1 -165 675 -165 675 7 Ibias
port 1 w
rlabel poly -165 645 -165 645 7 Vg
port 2 w
rlabel metal1 -165 300 -165 300 7 GND
port 3 w
rlabel locali -165 -780 -165 -780 7 Iout
port 4 w
rlabel poly 105 -835 105 -835 5 D0
port 5 s
rlabel poly 205 -835 205 -835 5 D0b
port 6 s
rlabel poly 805 -835 805 -835 5 D1
port 7 s
rlabel poly 905 -835 905 -835 5 D1b
port 8 s
rlabel poly 1505 -835 1505 -835 5 D2
port 9 s
rlabel poly 1605 -835 1605 -835 5 D2b
port 10 s
rlabel poly 2205 -835 2205 -835 5 D3
port 11 s
rlabel poly 2305 -835 2305 -835 5 D3b
port 12 s
rlabel poly 2905 -835 2905 -835 5 D4
port 13 s
rlabel poly 3005 -835 3005 -835 5 D4b
port 14 s
rlabel poly 3605 -835 3605 -835 5 D5
port 15 s
rlabel poly 3705 -835 3705 -835 5 D5b
port 16 s
rlabel poly 4305 -835 4305 -835 5 D6
port 17 s
rlabel poly 4405 -835 4405 -835 5 D6b
port 18 s
<< end >>

magic
tech sky130A
timestamp 1699199936
<< nwell >>
rect 690 850 1030 1675
rect 1390 850 1730 1675
rect 2090 850 2430 1675
rect 2790 850 3130 1675
rect 3490 850 3830 1675
rect 4190 850 4530 1675
<< nmos >>
rect 760 675 775 775
rect 800 675 815 775
rect 865 675 895 775
rect 945 675 960 775
rect 1460 675 1475 775
rect 1500 675 1515 775
rect 1565 675 1595 775
rect 1645 675 1660 775
rect 2160 675 2175 775
rect 2200 675 2215 775
rect 2265 675 2295 775
rect 2345 675 2360 775
rect 2860 675 2875 775
rect 2900 675 2915 775
rect 2965 675 2995 775
rect 3045 675 3060 775
rect 3560 675 3575 775
rect 3600 675 3615 775
rect 3665 675 3695 775
rect 3745 675 3760 775
rect 4260 675 4275 775
rect 4300 675 4315 775
rect 4365 675 4395 775
rect 4445 675 4460 775
rect 760 185 775 285
rect 800 185 815 285
rect 865 185 895 285
rect 945 185 960 285
rect 1460 185 1475 285
rect 1500 185 1515 285
rect 1565 185 1595 285
rect 1645 185 1660 285
rect 2160 185 2175 285
rect 2200 185 2215 285
rect 2265 185 2295 285
rect 2345 185 2360 285
rect 2860 185 2875 285
rect 2900 185 2915 285
rect 2965 185 2995 285
rect 3045 185 3060 285
rect 3560 185 3575 285
rect 3600 185 3615 285
rect 3665 185 3695 285
rect 3745 185 3760 285
rect 4260 185 4275 285
rect 4300 185 4315 285
rect 4365 185 4395 285
rect 4445 185 4460 285
<< pmos >>
rect 760 1400 775 1500
rect 825 1400 840 1500
rect 890 1400 905 1500
rect 945 1400 960 1500
rect 1460 1400 1475 1500
rect 1525 1400 1540 1500
rect 1590 1400 1605 1500
rect 1645 1400 1660 1500
rect 2160 1400 2175 1500
rect 2225 1400 2240 1500
rect 2290 1400 2305 1500
rect 2345 1400 2360 1500
rect 2860 1400 2875 1500
rect 2925 1400 2940 1500
rect 2990 1400 3005 1500
rect 3045 1400 3060 1500
rect 3560 1400 3575 1500
rect 3625 1400 3640 1500
rect 3690 1400 3705 1500
rect 3745 1400 3760 1500
rect 4260 1400 4275 1500
rect 4325 1400 4340 1500
rect 4390 1400 4405 1500
rect 4445 1400 4460 1500
rect 760 870 775 970
rect 825 870 840 970
rect 890 870 905 970
rect 945 870 960 970
rect 1460 870 1475 970
rect 1525 870 1540 970
rect 1590 870 1605 970
rect 1645 870 1660 970
rect 2160 870 2175 970
rect 2225 870 2240 970
rect 2290 870 2305 970
rect 2345 870 2360 970
rect 2860 870 2875 970
rect 2925 870 2940 970
rect 2990 870 3005 970
rect 3045 870 3060 970
rect 3560 870 3575 970
rect 3625 870 3640 970
rect 3690 870 3705 970
rect 3745 870 3760 970
rect 4260 870 4275 970
rect 4325 870 4340 970
rect 4390 870 4405 970
rect 4445 870 4460 970
<< ndiff >>
rect 710 760 760 775
rect 710 690 725 760
rect 745 690 760 760
rect 710 675 760 690
rect 775 675 800 775
rect 815 760 865 775
rect 815 690 830 760
rect 850 690 865 760
rect 815 675 865 690
rect 895 760 945 775
rect 895 690 910 760
rect 930 690 945 760
rect 895 675 945 690
rect 960 760 1010 775
rect 960 690 975 760
rect 995 690 1010 760
rect 960 675 1010 690
rect 1410 760 1460 775
rect 1410 690 1425 760
rect 1445 690 1460 760
rect 1410 675 1460 690
rect 1475 675 1500 775
rect 1515 760 1565 775
rect 1515 690 1530 760
rect 1550 690 1565 760
rect 1515 675 1565 690
rect 1595 760 1645 775
rect 1595 690 1610 760
rect 1630 690 1645 760
rect 1595 675 1645 690
rect 1660 760 1710 775
rect 1660 690 1675 760
rect 1695 690 1710 760
rect 1660 675 1710 690
rect 2110 760 2160 775
rect 2110 690 2125 760
rect 2145 690 2160 760
rect 2110 675 2160 690
rect 2175 675 2200 775
rect 2215 760 2265 775
rect 2215 690 2230 760
rect 2250 690 2265 760
rect 2215 675 2265 690
rect 2295 760 2345 775
rect 2295 690 2310 760
rect 2330 690 2345 760
rect 2295 675 2345 690
rect 2360 760 2410 775
rect 2360 690 2375 760
rect 2395 690 2410 760
rect 2360 675 2410 690
rect 2810 760 2860 775
rect 2810 690 2825 760
rect 2845 690 2860 760
rect 2810 675 2860 690
rect 2875 675 2900 775
rect 2915 760 2965 775
rect 2915 690 2930 760
rect 2950 690 2965 760
rect 2915 675 2965 690
rect 2995 760 3045 775
rect 2995 690 3010 760
rect 3030 690 3045 760
rect 2995 675 3045 690
rect 3060 760 3110 775
rect 3060 690 3075 760
rect 3095 690 3110 760
rect 3060 675 3110 690
rect 3510 760 3560 775
rect 3510 690 3525 760
rect 3545 690 3560 760
rect 3510 675 3560 690
rect 3575 675 3600 775
rect 3615 760 3665 775
rect 3615 690 3630 760
rect 3650 690 3665 760
rect 3615 675 3665 690
rect 3695 760 3745 775
rect 3695 690 3710 760
rect 3730 690 3745 760
rect 3695 675 3745 690
rect 3760 760 3810 775
rect 3760 690 3775 760
rect 3795 690 3810 760
rect 3760 675 3810 690
rect 4210 760 4260 775
rect 4210 690 4225 760
rect 4245 690 4260 760
rect 4210 675 4260 690
rect 4275 675 4300 775
rect 4315 760 4365 775
rect 4315 690 4330 760
rect 4350 690 4365 760
rect 4315 675 4365 690
rect 4395 760 4445 775
rect 4395 690 4410 760
rect 4430 690 4445 760
rect 4395 675 4445 690
rect 4460 760 4510 775
rect 4460 690 4475 760
rect 4495 690 4510 760
rect 4460 675 4510 690
rect 710 270 760 285
rect 710 200 725 270
rect 745 200 760 270
rect 710 185 760 200
rect 775 185 800 285
rect 815 270 865 285
rect 815 200 830 270
rect 850 200 865 270
rect 815 185 865 200
rect 895 270 945 285
rect 895 200 910 270
rect 930 200 945 270
rect 895 185 945 200
rect 960 270 1010 285
rect 960 200 975 270
rect 995 200 1010 270
rect 960 185 1010 200
rect 1410 270 1460 285
rect 1410 200 1425 270
rect 1445 200 1460 270
rect 1410 185 1460 200
rect 1475 185 1500 285
rect 1515 270 1565 285
rect 1515 200 1530 270
rect 1550 200 1565 270
rect 1515 185 1565 200
rect 1595 270 1645 285
rect 1595 200 1610 270
rect 1630 200 1645 270
rect 1595 185 1645 200
rect 1660 270 1710 285
rect 1660 200 1675 270
rect 1695 200 1710 270
rect 1660 185 1710 200
rect 2110 270 2160 285
rect 2110 200 2125 270
rect 2145 200 2160 270
rect 2110 185 2160 200
rect 2175 185 2200 285
rect 2215 270 2265 285
rect 2215 200 2230 270
rect 2250 200 2265 270
rect 2215 185 2265 200
rect 2295 270 2345 285
rect 2295 200 2310 270
rect 2330 200 2345 270
rect 2295 185 2345 200
rect 2360 270 2410 285
rect 2360 200 2375 270
rect 2395 200 2410 270
rect 2360 185 2410 200
rect 2810 270 2860 285
rect 2810 200 2825 270
rect 2845 200 2860 270
rect 2810 185 2860 200
rect 2875 185 2900 285
rect 2915 270 2965 285
rect 2915 200 2930 270
rect 2950 200 2965 270
rect 2915 185 2965 200
rect 2995 270 3045 285
rect 2995 200 3010 270
rect 3030 200 3045 270
rect 2995 185 3045 200
rect 3060 270 3110 285
rect 3060 200 3075 270
rect 3095 200 3110 270
rect 3060 185 3110 200
rect 3510 270 3560 285
rect 3510 200 3525 270
rect 3545 200 3560 270
rect 3510 185 3560 200
rect 3575 185 3600 285
rect 3615 270 3665 285
rect 3615 200 3630 270
rect 3650 200 3665 270
rect 3615 185 3665 200
rect 3695 270 3745 285
rect 3695 200 3710 270
rect 3730 200 3745 270
rect 3695 185 3745 200
rect 3760 270 3810 285
rect 3760 200 3775 270
rect 3795 200 3810 270
rect 3760 185 3810 200
rect 4210 270 4260 285
rect 4210 200 4225 270
rect 4245 200 4260 270
rect 4210 185 4260 200
rect 4275 185 4300 285
rect 4315 270 4365 285
rect 4315 200 4330 270
rect 4350 200 4365 270
rect 4315 185 4365 200
rect 4395 270 4445 285
rect 4395 200 4410 270
rect 4430 200 4445 270
rect 4395 185 4445 200
rect 4460 270 4510 285
rect 4460 200 4475 270
rect 4495 200 4510 270
rect 4460 185 4510 200
<< pdiff >>
rect 710 1485 760 1500
rect 710 1415 725 1485
rect 745 1415 760 1485
rect 710 1400 760 1415
rect 775 1485 825 1500
rect 775 1415 790 1485
rect 810 1415 825 1485
rect 775 1400 825 1415
rect 840 1485 890 1500
rect 840 1415 855 1485
rect 875 1415 890 1485
rect 840 1400 890 1415
rect 905 1400 945 1500
rect 960 1485 1010 1500
rect 960 1415 975 1485
rect 995 1415 1010 1485
rect 960 1400 1010 1415
rect 1410 1485 1460 1500
rect 1410 1415 1425 1485
rect 1445 1415 1460 1485
rect 1410 1400 1460 1415
rect 1475 1485 1525 1500
rect 1475 1415 1490 1485
rect 1510 1415 1525 1485
rect 1475 1400 1525 1415
rect 1540 1485 1590 1500
rect 1540 1415 1555 1485
rect 1575 1415 1590 1485
rect 1540 1400 1590 1415
rect 1605 1400 1645 1500
rect 1660 1485 1710 1500
rect 1660 1415 1675 1485
rect 1695 1415 1710 1485
rect 1660 1400 1710 1415
rect 2110 1485 2160 1500
rect 2110 1415 2125 1485
rect 2145 1415 2160 1485
rect 2110 1400 2160 1415
rect 2175 1485 2225 1500
rect 2175 1415 2190 1485
rect 2210 1415 2225 1485
rect 2175 1400 2225 1415
rect 2240 1485 2290 1500
rect 2240 1415 2255 1485
rect 2275 1415 2290 1485
rect 2240 1400 2290 1415
rect 2305 1400 2345 1500
rect 2360 1485 2410 1500
rect 2360 1415 2375 1485
rect 2395 1415 2410 1485
rect 2360 1400 2410 1415
rect 2810 1485 2860 1500
rect 2810 1415 2825 1485
rect 2845 1415 2860 1485
rect 2810 1400 2860 1415
rect 2875 1485 2925 1500
rect 2875 1415 2890 1485
rect 2910 1415 2925 1485
rect 2875 1400 2925 1415
rect 2940 1485 2990 1500
rect 2940 1415 2955 1485
rect 2975 1415 2990 1485
rect 2940 1400 2990 1415
rect 3005 1400 3045 1500
rect 3060 1485 3110 1500
rect 3060 1415 3075 1485
rect 3095 1415 3110 1485
rect 3060 1400 3110 1415
rect 3510 1485 3560 1500
rect 3510 1415 3525 1485
rect 3545 1415 3560 1485
rect 3510 1400 3560 1415
rect 3575 1485 3625 1500
rect 3575 1415 3590 1485
rect 3610 1415 3625 1485
rect 3575 1400 3625 1415
rect 3640 1485 3690 1500
rect 3640 1415 3655 1485
rect 3675 1415 3690 1485
rect 3640 1400 3690 1415
rect 3705 1400 3745 1500
rect 3760 1485 3810 1500
rect 3760 1415 3775 1485
rect 3795 1415 3810 1485
rect 3760 1400 3810 1415
rect 4210 1485 4260 1500
rect 4210 1415 4225 1485
rect 4245 1415 4260 1485
rect 4210 1400 4260 1415
rect 4275 1485 4325 1500
rect 4275 1415 4290 1485
rect 4310 1415 4325 1485
rect 4275 1400 4325 1415
rect 4340 1485 4390 1500
rect 4340 1415 4355 1485
rect 4375 1415 4390 1485
rect 4340 1400 4390 1415
rect 4405 1400 4445 1500
rect 4460 1485 4510 1500
rect 4460 1415 4475 1485
rect 4495 1415 4510 1485
rect 4460 1400 4510 1415
rect 710 955 760 970
rect 710 885 725 955
rect 745 885 760 955
rect 710 870 760 885
rect 775 955 825 970
rect 775 885 790 955
rect 810 885 825 955
rect 775 870 825 885
rect 840 955 890 970
rect 840 885 855 955
rect 875 885 890 955
rect 840 870 890 885
rect 905 870 945 970
rect 960 955 1010 970
rect 960 885 975 955
rect 995 885 1010 955
rect 960 870 1010 885
rect 1410 955 1460 970
rect 1410 885 1425 955
rect 1445 885 1460 955
rect 1410 870 1460 885
rect 1475 955 1525 970
rect 1475 885 1490 955
rect 1510 885 1525 955
rect 1475 870 1525 885
rect 1540 955 1590 970
rect 1540 885 1555 955
rect 1575 885 1590 955
rect 1540 870 1590 885
rect 1605 870 1645 970
rect 1660 955 1710 970
rect 1660 885 1675 955
rect 1695 885 1710 955
rect 1660 870 1710 885
rect 2110 955 2160 970
rect 2110 885 2125 955
rect 2145 885 2160 955
rect 2110 870 2160 885
rect 2175 955 2225 970
rect 2175 885 2190 955
rect 2210 885 2225 955
rect 2175 870 2225 885
rect 2240 955 2290 970
rect 2240 885 2255 955
rect 2275 885 2290 955
rect 2240 870 2290 885
rect 2305 870 2345 970
rect 2360 955 2410 970
rect 2360 885 2375 955
rect 2395 885 2410 955
rect 2360 870 2410 885
rect 2810 955 2860 970
rect 2810 885 2825 955
rect 2845 885 2860 955
rect 2810 870 2860 885
rect 2875 955 2925 970
rect 2875 885 2890 955
rect 2910 885 2925 955
rect 2875 870 2925 885
rect 2940 955 2990 970
rect 2940 885 2955 955
rect 2975 885 2990 955
rect 2940 870 2990 885
rect 3005 870 3045 970
rect 3060 955 3110 970
rect 3060 885 3075 955
rect 3095 885 3110 955
rect 3060 870 3110 885
rect 3510 955 3560 970
rect 3510 885 3525 955
rect 3545 885 3560 955
rect 3510 870 3560 885
rect 3575 955 3625 970
rect 3575 885 3590 955
rect 3610 885 3625 955
rect 3575 870 3625 885
rect 3640 955 3690 970
rect 3640 885 3655 955
rect 3675 885 3690 955
rect 3640 870 3690 885
rect 3705 870 3745 970
rect 3760 955 3810 970
rect 3760 885 3775 955
rect 3795 885 3810 955
rect 3760 870 3810 885
rect 4210 955 4260 970
rect 4210 885 4225 955
rect 4245 885 4260 955
rect 4210 870 4260 885
rect 4275 955 4325 970
rect 4275 885 4290 955
rect 4310 885 4325 955
rect 4275 870 4325 885
rect 4340 955 4390 970
rect 4340 885 4355 955
rect 4375 885 4390 955
rect 4340 870 4390 885
rect 4405 870 4445 970
rect 4460 955 4510 970
rect 4460 885 4475 955
rect 4495 885 4510 955
rect 4460 870 4510 885
<< ndiffc >>
rect 725 690 745 760
rect 830 690 850 760
rect 910 690 930 760
rect 975 690 995 760
rect 1425 690 1445 760
rect 1530 690 1550 760
rect 1610 690 1630 760
rect 1675 690 1695 760
rect 2125 690 2145 760
rect 2230 690 2250 760
rect 2310 690 2330 760
rect 2375 690 2395 760
rect 2825 690 2845 760
rect 2930 690 2950 760
rect 3010 690 3030 760
rect 3075 690 3095 760
rect 3525 690 3545 760
rect 3630 690 3650 760
rect 3710 690 3730 760
rect 3775 690 3795 760
rect 4225 690 4245 760
rect 4330 690 4350 760
rect 4410 690 4430 760
rect 4475 690 4495 760
rect 725 200 745 270
rect 830 200 850 270
rect 910 200 930 270
rect 975 200 995 270
rect 1425 200 1445 270
rect 1530 200 1550 270
rect 1610 200 1630 270
rect 1675 200 1695 270
rect 2125 200 2145 270
rect 2230 200 2250 270
rect 2310 200 2330 270
rect 2375 200 2395 270
rect 2825 200 2845 270
rect 2930 200 2950 270
rect 3010 200 3030 270
rect 3075 200 3095 270
rect 3525 200 3545 270
rect 3630 200 3650 270
rect 3710 200 3730 270
rect 3775 200 3795 270
rect 4225 200 4245 270
rect 4330 200 4350 270
rect 4410 200 4430 270
rect 4475 200 4495 270
<< pdiffc >>
rect 725 1415 745 1485
rect 790 1415 810 1485
rect 855 1415 875 1485
rect 975 1415 995 1485
rect 1425 1415 1445 1485
rect 1490 1415 1510 1485
rect 1555 1415 1575 1485
rect 1675 1415 1695 1485
rect 2125 1415 2145 1485
rect 2190 1415 2210 1485
rect 2255 1415 2275 1485
rect 2375 1415 2395 1485
rect 2825 1415 2845 1485
rect 2890 1415 2910 1485
rect 2955 1415 2975 1485
rect 3075 1415 3095 1485
rect 3525 1415 3545 1485
rect 3590 1415 3610 1485
rect 3655 1415 3675 1485
rect 3775 1415 3795 1485
rect 4225 1415 4245 1485
rect 4290 1415 4310 1485
rect 4355 1415 4375 1485
rect 4475 1415 4495 1485
rect 725 885 745 955
rect 790 885 810 955
rect 855 885 875 955
rect 975 885 995 955
rect 1425 885 1445 955
rect 1490 885 1510 955
rect 1555 885 1575 955
rect 1675 885 1695 955
rect 2125 885 2145 955
rect 2190 885 2210 955
rect 2255 885 2275 955
rect 2375 885 2395 955
rect 2825 885 2845 955
rect 2890 885 2910 955
rect 2955 885 2975 955
rect 3075 885 3095 955
rect 3525 885 3545 955
rect 3590 885 3610 955
rect 3655 885 3675 955
rect 3775 885 3795 955
rect 4225 885 4245 955
rect 4290 885 4310 955
rect 4355 885 4375 955
rect 4475 885 4495 955
<< psubdiff >>
rect 785 140 835 155
rect 785 70 800 140
rect 820 70 835 140
rect 785 55 835 70
rect 920 140 970 155
rect 920 70 935 140
rect 955 70 970 140
rect 920 55 970 70
rect 1485 140 1535 155
rect 1485 70 1500 140
rect 1520 70 1535 140
rect 1485 55 1535 70
rect 1620 140 1670 155
rect 1620 70 1635 140
rect 1655 70 1670 140
rect 1620 55 1670 70
rect 2185 140 2235 155
rect 2185 70 2200 140
rect 2220 70 2235 140
rect 2185 55 2235 70
rect 2320 140 2370 155
rect 2320 70 2335 140
rect 2355 70 2370 140
rect 2320 55 2370 70
rect 2885 140 2935 155
rect 2885 70 2900 140
rect 2920 70 2935 140
rect 2885 55 2935 70
rect 3020 140 3070 155
rect 3020 70 3035 140
rect 3055 70 3070 140
rect 3020 55 3070 70
rect 3585 140 3635 155
rect 3585 70 3600 140
rect 3620 70 3635 140
rect 3585 55 3635 70
rect 3720 140 3770 155
rect 3720 70 3735 140
rect 3755 70 3770 140
rect 3720 55 3770 70
rect 4285 140 4335 155
rect 4285 70 4300 140
rect 4320 70 4335 140
rect 4285 55 4335 70
rect 4420 140 4470 155
rect 4420 70 4435 140
rect 4455 70 4470 140
rect 4420 55 4470 70
<< nsubdiff >>
rect 765 1640 815 1655
rect 765 1570 780 1640
rect 800 1570 815 1640
rect 765 1555 815 1570
rect 905 1640 955 1655
rect 905 1570 920 1640
rect 940 1570 955 1640
rect 1465 1640 1515 1655
rect 905 1555 955 1570
rect 1465 1570 1480 1640
rect 1500 1570 1515 1640
rect 1465 1555 1515 1570
rect 1605 1640 1655 1655
rect 1605 1570 1620 1640
rect 1640 1570 1655 1640
rect 2165 1640 2215 1655
rect 1605 1555 1655 1570
rect 2165 1570 2180 1640
rect 2200 1570 2215 1640
rect 2165 1555 2215 1570
rect 2305 1640 2355 1655
rect 2305 1570 2320 1640
rect 2340 1570 2355 1640
rect 2865 1640 2915 1655
rect 2305 1555 2355 1570
rect 2865 1570 2880 1640
rect 2900 1570 2915 1640
rect 2865 1555 2915 1570
rect 3005 1640 3055 1655
rect 3005 1570 3020 1640
rect 3040 1570 3055 1640
rect 3565 1640 3615 1655
rect 3005 1555 3055 1570
rect 3565 1570 3580 1640
rect 3600 1570 3615 1640
rect 3565 1555 3615 1570
rect 3705 1640 3755 1655
rect 3705 1570 3720 1640
rect 3740 1570 3755 1640
rect 4265 1640 4315 1655
rect 3705 1555 3755 1570
rect 4265 1570 4280 1640
rect 4300 1570 4315 1640
rect 4265 1555 4315 1570
rect 4405 1640 4455 1655
rect 4405 1570 4420 1640
rect 4440 1570 4455 1640
rect 4405 1555 4455 1570
<< psubdiffcont >>
rect 800 70 820 140
rect 935 70 955 140
rect 1500 70 1520 140
rect 1635 70 1655 140
rect 2200 70 2220 140
rect 2335 70 2355 140
rect 2900 70 2920 140
rect 3035 70 3055 140
rect 3600 70 3620 140
rect 3735 70 3755 140
rect 4300 70 4320 140
rect 4435 70 4455 140
<< nsubdiffcont >>
rect 780 1570 800 1640
rect 920 1570 940 1640
rect 1480 1570 1500 1640
rect 1620 1570 1640 1640
rect 2180 1570 2200 1640
rect 2320 1570 2340 1640
rect 2880 1570 2900 1640
rect 3020 1570 3040 1640
rect 3580 1570 3600 1640
rect 3720 1570 3740 1640
rect 4280 1570 4300 1640
rect 4420 1570 4440 1640
<< poly >>
rect 1655 1700 1670 1710
rect 270 1670 285 1700
rect 355 1670 370 1685
rect 970 1670 985 1695
rect 1055 1670 1070 1685
rect 1655 1680 1685 1700
rect 1670 1670 1685 1680
rect 1755 1670 1770 1710
rect 2355 1695 2370 1710
rect 2355 1680 2385 1695
rect 2370 1670 2385 1680
rect 2455 1670 2470 1710
rect 3055 1700 3070 1710
rect 3055 1680 3085 1700
rect 3070 1670 3085 1680
rect 3155 1670 3170 1710
rect 3755 1695 3770 1710
rect 3755 1680 3785 1695
rect 3770 1670 3785 1680
rect 3855 1670 3870 1710
rect 4455 1700 4470 1710
rect 4455 1680 4485 1700
rect 4470 1670 4485 1680
rect 4555 1670 4570 1710
rect 270 1660 310 1670
rect 270 1640 280 1660
rect 300 1640 310 1660
rect 270 1630 310 1640
rect 335 1660 375 1670
rect 335 1640 345 1660
rect 365 1640 375 1660
rect 970 1660 1010 1670
rect 335 1630 375 1640
rect 970 1640 980 1660
rect 1000 1640 1010 1660
rect 970 1630 1010 1640
rect 1035 1660 1075 1670
rect 1035 1640 1045 1660
rect 1065 1640 1075 1660
rect 1670 1660 1710 1670
rect 1035 1630 1075 1640
rect 1670 1640 1680 1660
rect 1700 1640 1710 1660
rect 1670 1630 1710 1640
rect 1735 1660 1775 1670
rect 1735 1640 1745 1660
rect 1765 1640 1775 1660
rect 2370 1660 2410 1670
rect 1735 1630 1775 1640
rect 2370 1640 2380 1660
rect 2400 1640 2410 1660
rect 2370 1630 2410 1640
rect 2435 1660 2475 1670
rect 2435 1640 2445 1660
rect 2465 1640 2475 1660
rect 3070 1660 3110 1670
rect 2435 1630 2475 1640
rect 3070 1640 3080 1660
rect 3100 1640 3110 1660
rect 3070 1630 3110 1640
rect 3135 1660 3175 1670
rect 3135 1640 3145 1660
rect 3165 1640 3175 1660
rect 3770 1660 3810 1670
rect 3135 1630 3175 1640
rect 3770 1640 3780 1660
rect 3800 1640 3810 1660
rect 3770 1630 3810 1640
rect 3835 1660 3875 1670
rect 3835 1640 3845 1660
rect 3865 1640 3875 1660
rect 4470 1660 4510 1670
rect 3835 1630 3875 1640
rect 4470 1640 4480 1660
rect 4500 1640 4510 1660
rect 4470 1630 4510 1640
rect 4535 1660 4575 1670
rect 4535 1640 4545 1660
rect 4565 1640 4575 1660
rect 4535 1630 4575 1640
rect 760 1500 775 1515
rect 825 1500 840 1515
rect 890 1500 905 1515
rect 945 1500 960 1515
rect 1460 1500 1475 1515
rect 1525 1500 1540 1515
rect 1590 1500 1605 1515
rect 1645 1500 1660 1515
rect 2160 1500 2175 1515
rect 2225 1500 2240 1515
rect 2290 1500 2305 1515
rect 2345 1500 2360 1515
rect 2860 1500 2875 1515
rect 2925 1500 2940 1515
rect 2990 1500 3005 1515
rect 3045 1500 3060 1515
rect 3560 1500 3575 1515
rect 3625 1500 3640 1515
rect 3690 1500 3705 1515
rect 3745 1500 3760 1515
rect 4260 1500 4275 1515
rect 4325 1500 4340 1515
rect 4390 1500 4405 1515
rect 4445 1500 4460 1515
rect 760 1365 775 1400
rect 760 1350 800 1365
rect 785 1175 800 1350
rect 760 1160 800 1175
rect 760 970 775 1160
rect 825 1135 840 1400
rect 800 1125 840 1135
rect 800 1105 810 1125
rect 830 1105 840 1125
rect 800 1095 840 1105
rect 800 1060 840 1070
rect 800 1040 810 1060
rect 830 1040 840 1060
rect 800 1030 840 1040
rect 825 970 840 1030
rect 890 970 905 1400
rect 945 1340 960 1400
rect 1460 1365 1475 1400
rect 1460 1350 1500 1365
rect 930 1330 970 1340
rect 930 1310 940 1330
rect 960 1310 970 1330
rect 930 1300 970 1310
rect 930 1265 970 1275
rect 930 1245 940 1265
rect 960 1245 970 1265
rect 930 1235 970 1245
rect 945 970 960 1235
rect 1485 1175 1500 1350
rect 1460 1160 1500 1175
rect 1460 970 1475 1160
rect 1525 1135 1540 1400
rect 1500 1125 1540 1135
rect 1500 1105 1510 1125
rect 1530 1105 1540 1125
rect 1500 1095 1540 1105
rect 1500 1060 1540 1070
rect 1500 1040 1510 1060
rect 1530 1040 1540 1060
rect 1500 1030 1540 1040
rect 1525 970 1540 1030
rect 1590 970 1605 1400
rect 1645 1340 1660 1400
rect 2160 1365 2175 1400
rect 2160 1350 2200 1365
rect 1630 1330 1670 1340
rect 1630 1310 1640 1330
rect 1660 1310 1670 1330
rect 1630 1300 1670 1310
rect 1630 1265 1670 1275
rect 1630 1245 1640 1265
rect 1660 1245 1670 1265
rect 1630 1235 1670 1245
rect 1645 970 1660 1235
rect 2185 1175 2200 1350
rect 2160 1160 2200 1175
rect 2160 970 2175 1160
rect 2225 1135 2240 1400
rect 2200 1125 2240 1135
rect 2200 1105 2210 1125
rect 2230 1105 2240 1125
rect 2200 1095 2240 1105
rect 2200 1060 2240 1070
rect 2200 1040 2210 1060
rect 2230 1040 2240 1060
rect 2200 1030 2240 1040
rect 2225 970 2240 1030
rect 2290 970 2305 1400
rect 2345 1340 2360 1400
rect 2860 1365 2875 1400
rect 2860 1350 2900 1365
rect 2330 1330 2370 1340
rect 2330 1310 2340 1330
rect 2360 1310 2370 1330
rect 2330 1300 2370 1310
rect 2330 1265 2370 1275
rect 2330 1245 2340 1265
rect 2360 1245 2370 1265
rect 2330 1235 2370 1245
rect 2345 970 2360 1235
rect 2885 1175 2900 1350
rect 2860 1160 2900 1175
rect 2860 970 2875 1160
rect 2925 1135 2940 1400
rect 2900 1125 2940 1135
rect 2900 1105 2910 1125
rect 2930 1105 2940 1125
rect 2900 1095 2940 1105
rect 2900 1060 2940 1070
rect 2900 1040 2910 1060
rect 2930 1040 2940 1060
rect 2900 1030 2940 1040
rect 2925 970 2940 1030
rect 2990 970 3005 1400
rect 3045 1340 3060 1400
rect 3560 1365 3575 1400
rect 3560 1350 3600 1365
rect 3030 1330 3070 1340
rect 3030 1310 3040 1330
rect 3060 1310 3070 1330
rect 3030 1300 3070 1310
rect 3030 1265 3070 1275
rect 3030 1245 3040 1265
rect 3060 1245 3070 1265
rect 3030 1235 3070 1245
rect 3045 970 3060 1235
rect 3585 1175 3600 1350
rect 3560 1160 3600 1175
rect 3560 970 3575 1160
rect 3625 1135 3640 1400
rect 3600 1125 3640 1135
rect 3600 1105 3610 1125
rect 3630 1105 3640 1125
rect 3600 1095 3640 1105
rect 3600 1060 3640 1070
rect 3600 1040 3610 1060
rect 3630 1040 3640 1060
rect 3600 1030 3640 1040
rect 3625 970 3640 1030
rect 3690 970 3705 1400
rect 3745 1340 3760 1400
rect 4260 1365 4275 1400
rect 4260 1350 4300 1365
rect 3730 1330 3770 1340
rect 3730 1310 3740 1330
rect 3760 1310 3770 1330
rect 3730 1300 3770 1310
rect 3730 1265 3770 1275
rect 3730 1245 3740 1265
rect 3760 1245 3770 1265
rect 3730 1235 3770 1245
rect 3745 970 3760 1235
rect 4285 1175 4300 1350
rect 4260 1160 4300 1175
rect 4260 970 4275 1160
rect 4325 1135 4340 1400
rect 4300 1125 4340 1135
rect 4300 1105 4310 1125
rect 4330 1105 4340 1125
rect 4300 1095 4340 1105
rect 4300 1060 4340 1070
rect 4300 1040 4310 1060
rect 4330 1040 4340 1060
rect 4300 1030 4340 1040
rect 4325 970 4340 1030
rect 4390 970 4405 1400
rect 4445 1340 4460 1400
rect 4430 1330 4470 1340
rect 4430 1310 4440 1330
rect 4460 1310 4470 1330
rect 4430 1300 4470 1310
rect 4430 1265 4470 1275
rect 4430 1245 4440 1265
rect 4460 1245 4470 1265
rect 4430 1235 4470 1245
rect 4445 970 4460 1235
rect 760 775 775 870
rect 825 855 840 870
rect 890 855 905 870
rect 800 840 840 855
rect 880 840 905 855
rect 800 775 815 840
rect 880 790 895 840
rect 865 775 895 790
rect 945 775 960 870
rect 1460 775 1475 870
rect 1525 855 1540 870
rect 1590 855 1605 870
rect 1500 840 1540 855
rect 1580 840 1605 855
rect 1500 775 1515 840
rect 1580 790 1595 840
rect 1565 775 1595 790
rect 1645 775 1660 870
rect 2160 775 2175 870
rect 2225 855 2240 870
rect 2290 855 2305 870
rect 2200 840 2240 855
rect 2280 840 2305 855
rect 2200 775 2215 840
rect 2280 790 2295 840
rect 2265 775 2295 790
rect 2345 775 2360 870
rect 2860 775 2875 870
rect 2925 855 2940 870
rect 2990 855 3005 870
rect 2900 840 2940 855
rect 2980 840 3005 855
rect 2900 775 2915 840
rect 2980 790 2995 840
rect 2965 775 2995 790
rect 3045 775 3060 870
rect 3560 775 3575 870
rect 3625 855 3640 870
rect 3690 855 3705 870
rect 3600 840 3640 855
rect 3680 840 3705 855
rect 3600 775 3615 840
rect 3680 790 3695 840
rect 3665 775 3695 790
rect 3745 775 3760 870
rect 4260 775 4275 870
rect 4325 855 4340 870
rect 4390 855 4405 870
rect 4300 840 4340 855
rect 4380 840 4405 855
rect 4300 775 4315 840
rect 4380 790 4395 840
rect 4365 775 4395 790
rect 4445 775 4460 870
rect 760 490 775 675
rect 800 620 815 675
rect 800 610 840 620
rect 800 590 810 610
rect 830 590 840 610
rect 800 580 840 590
rect 800 545 840 555
rect 800 525 810 545
rect 830 525 840 545
rect 800 515 840 525
rect 760 475 800 490
rect 785 355 800 475
rect 760 340 800 355
rect 760 285 775 340
rect 825 315 840 515
rect 800 300 840 315
rect 800 285 815 300
rect 865 285 895 675
rect 945 510 960 675
rect 945 495 980 510
rect 965 465 980 495
rect 1460 490 1475 675
rect 1500 620 1515 675
rect 1500 610 1540 620
rect 1500 590 1510 610
rect 1530 590 1540 610
rect 1500 580 1540 590
rect 1500 545 1540 555
rect 1500 525 1510 545
rect 1530 525 1540 545
rect 1500 515 1540 525
rect 1460 475 1500 490
rect 940 455 980 465
rect 940 435 950 455
rect 970 435 980 455
rect 940 425 980 435
rect 920 375 960 385
rect 920 355 930 375
rect 950 355 960 375
rect 1485 355 1500 475
rect 920 345 960 355
rect 945 285 960 345
rect 1460 340 1500 355
rect 1460 285 1475 340
rect 1525 315 1540 515
rect 1500 300 1540 315
rect 1500 285 1515 300
rect 1565 285 1595 675
rect 1645 510 1660 675
rect 1645 495 1680 510
rect 1665 465 1680 495
rect 2160 490 2175 675
rect 2200 620 2215 675
rect 2200 610 2240 620
rect 2200 590 2210 610
rect 2230 590 2240 610
rect 2200 580 2240 590
rect 2200 545 2240 555
rect 2200 525 2210 545
rect 2230 525 2240 545
rect 2200 515 2240 525
rect 2160 475 2200 490
rect 1640 455 1680 465
rect 1640 435 1650 455
rect 1670 435 1680 455
rect 1640 425 1680 435
rect 1620 375 1660 385
rect 1620 355 1630 375
rect 1650 355 1660 375
rect 2185 355 2200 475
rect 1620 345 1660 355
rect 1645 285 1660 345
rect 2160 340 2200 355
rect 2160 285 2175 340
rect 2225 315 2240 515
rect 2200 300 2240 315
rect 2200 285 2215 300
rect 2265 285 2295 675
rect 2345 510 2360 675
rect 2345 495 2380 510
rect 2365 465 2380 495
rect 2860 490 2875 675
rect 2900 620 2915 675
rect 2900 610 2940 620
rect 2900 590 2910 610
rect 2930 590 2940 610
rect 2900 580 2940 590
rect 2900 545 2940 555
rect 2900 525 2910 545
rect 2930 525 2940 545
rect 2900 515 2940 525
rect 2860 475 2900 490
rect 2340 455 2380 465
rect 2340 435 2350 455
rect 2370 435 2380 455
rect 2340 425 2380 435
rect 2320 375 2360 385
rect 2320 355 2330 375
rect 2350 355 2360 375
rect 2885 355 2900 475
rect 2320 345 2360 355
rect 2345 285 2360 345
rect 2860 340 2900 355
rect 2860 285 2875 340
rect 2925 315 2940 515
rect 2900 300 2940 315
rect 2900 285 2915 300
rect 2965 285 2995 675
rect 3045 510 3060 675
rect 3045 495 3080 510
rect 3065 465 3080 495
rect 3560 490 3575 675
rect 3600 620 3615 675
rect 3600 610 3640 620
rect 3600 590 3610 610
rect 3630 590 3640 610
rect 3600 580 3640 590
rect 3600 545 3640 555
rect 3600 525 3610 545
rect 3630 525 3640 545
rect 3600 515 3640 525
rect 3560 475 3600 490
rect 3040 455 3080 465
rect 3040 435 3050 455
rect 3070 435 3080 455
rect 3040 425 3080 435
rect 3020 375 3060 385
rect 3020 355 3030 375
rect 3050 355 3060 375
rect 3585 355 3600 475
rect 3020 345 3060 355
rect 3045 285 3060 345
rect 3560 340 3600 355
rect 3560 285 3575 340
rect 3625 315 3640 515
rect 3600 300 3640 315
rect 3600 285 3615 300
rect 3665 285 3695 675
rect 3745 510 3760 675
rect 3745 495 3780 510
rect 3765 465 3780 495
rect 4260 490 4275 675
rect 4300 620 4315 675
rect 4300 610 4340 620
rect 4300 590 4310 610
rect 4330 590 4340 610
rect 4300 580 4340 590
rect 4300 545 4340 555
rect 4300 525 4310 545
rect 4330 525 4340 545
rect 4300 515 4340 525
rect 4260 475 4300 490
rect 3740 455 3780 465
rect 3740 435 3750 455
rect 3770 435 3780 455
rect 3740 425 3780 435
rect 3720 375 3760 385
rect 3720 355 3730 375
rect 3750 355 3760 375
rect 4285 355 4300 475
rect 3720 345 3760 355
rect 3745 285 3760 345
rect 4260 340 4300 355
rect 4260 285 4275 340
rect 4325 315 4340 515
rect 4300 300 4340 315
rect 4300 285 4315 300
rect 4365 285 4395 675
rect 4445 510 4460 675
rect 4445 495 4480 510
rect 4465 465 4480 495
rect 4440 455 4480 465
rect 4440 435 4450 455
rect 4470 435 4480 455
rect 4440 425 4480 435
rect 4420 375 4460 385
rect 4420 355 4430 375
rect 4450 355 4460 375
rect 4420 345 4460 355
rect 4445 285 4460 345
rect 760 40 775 185
rect 800 170 815 185
rect 865 40 895 185
rect 945 170 960 185
rect 1460 40 1475 185
rect 1500 170 1515 185
rect 1565 40 1595 185
rect 1645 170 1660 185
rect 2160 40 2175 185
rect 2200 170 2215 185
rect 2265 40 2295 185
rect 2345 170 2360 185
rect 2860 40 2875 185
rect 2900 170 2915 185
rect 2965 40 2995 185
rect 3045 170 3060 185
rect 3560 40 3575 185
rect 3600 170 3615 185
rect 3665 40 3695 185
rect 3745 170 3760 185
rect 4260 40 4275 185
rect 4300 170 4315 185
rect 4365 40 4395 185
rect 4445 170 4460 185
rect 735 30 775 40
rect 735 10 745 30
rect 765 10 775 30
rect 735 0 775 10
rect 855 30 895 40
rect 855 10 865 30
rect 885 10 895 30
rect 855 0 895 10
rect 1435 30 1475 40
rect 1435 10 1445 30
rect 1465 10 1475 30
rect 1435 0 1475 10
rect 1555 30 1595 40
rect 1555 10 1565 30
rect 1585 10 1595 30
rect 1555 0 1595 10
rect 2135 30 2175 40
rect 2135 10 2145 30
rect 2165 10 2175 30
rect 2135 0 2175 10
rect 2255 30 2295 40
rect 2255 10 2265 30
rect 2285 10 2295 30
rect 2255 0 2295 10
rect 2835 30 2875 40
rect 2835 10 2845 30
rect 2865 10 2875 30
rect 2835 0 2875 10
rect 2955 30 2995 40
rect 2955 10 2965 30
rect 2985 10 2995 30
rect 2955 0 2995 10
rect 3535 30 3575 40
rect 3535 10 3545 30
rect 3565 10 3575 30
rect 3535 0 3575 10
rect 3655 30 3695 40
rect 3655 10 3665 30
rect 3685 10 3695 30
rect 3655 0 3695 10
rect 4235 30 4275 40
rect 4235 10 4245 30
rect 4265 10 4275 30
rect 4235 0 4275 10
rect 4355 30 4395 40
rect 4355 10 4365 30
rect 4385 10 4395 30
rect 4355 0 4395 10
<< polycont >>
rect 280 1640 300 1660
rect 345 1640 365 1660
rect 980 1640 1000 1660
rect 1045 1640 1065 1660
rect 1680 1640 1700 1660
rect 1745 1640 1765 1660
rect 2380 1640 2400 1660
rect 2445 1640 2465 1660
rect 3080 1640 3100 1660
rect 3145 1640 3165 1660
rect 3780 1640 3800 1660
rect 3845 1640 3865 1660
rect 4480 1640 4500 1660
rect 4545 1640 4565 1660
rect 810 1105 830 1125
rect 810 1040 830 1060
rect 940 1310 960 1330
rect 940 1245 960 1265
rect 1510 1105 1530 1125
rect 1510 1040 1530 1060
rect 1640 1310 1660 1330
rect 1640 1245 1660 1265
rect 2210 1105 2230 1125
rect 2210 1040 2230 1060
rect 2340 1310 2360 1330
rect 2340 1245 2360 1265
rect 2910 1105 2930 1125
rect 2910 1040 2930 1060
rect 3040 1310 3060 1330
rect 3040 1245 3060 1265
rect 3610 1105 3630 1125
rect 3610 1040 3630 1060
rect 3740 1310 3760 1330
rect 3740 1245 3760 1265
rect 4310 1105 4330 1125
rect 4310 1040 4330 1060
rect 4440 1310 4460 1330
rect 4440 1245 4460 1265
rect 810 590 830 610
rect 810 525 830 545
rect 1510 590 1530 610
rect 1510 525 1530 545
rect 950 435 970 455
rect 930 355 950 375
rect 2210 590 2230 610
rect 2210 525 2230 545
rect 1650 435 1670 455
rect 1630 355 1650 375
rect 2910 590 2930 610
rect 2910 525 2930 545
rect 2350 435 2370 455
rect 2330 355 2350 375
rect 3610 590 3630 610
rect 3610 525 3630 545
rect 3050 435 3070 455
rect 3030 355 3050 375
rect 4310 590 4330 610
rect 4310 525 4330 545
rect 3750 435 3770 455
rect 3730 355 3750 375
rect 4450 435 4470 455
rect 4430 355 4450 375
rect 745 10 765 30
rect 865 10 885 30
rect 1445 10 1465 30
rect 1565 10 1585 30
rect 2145 10 2165 30
rect 2265 10 2285 30
rect 2845 10 2865 30
rect 2965 10 2985 30
rect 3545 10 3565 30
rect 3665 10 3685 30
rect 4245 10 4265 30
rect 4365 10 4385 30
<< locali >>
rect 270 1660 310 1670
rect 270 1640 280 1660
rect 300 1640 310 1660
rect 270 1630 310 1640
rect 335 1660 375 1670
rect 335 1640 345 1660
rect 365 1640 375 1660
rect 970 1660 1010 1670
rect 335 1630 375 1640
rect 770 1640 810 1650
rect 285 1495 305 1630
rect 335 965 355 1630
rect 770 1570 780 1640
rect 800 1570 810 1640
rect 770 1560 810 1570
rect 910 1640 950 1650
rect 910 1570 920 1640
rect 940 1570 950 1640
rect 970 1640 980 1660
rect 1000 1640 1010 1660
rect 970 1630 1010 1640
rect 1035 1660 1075 1670
rect 1035 1640 1045 1660
rect 1065 1640 1075 1660
rect 1670 1660 1710 1670
rect 1035 1630 1075 1640
rect 1470 1640 1510 1650
rect 910 1560 950 1570
rect 985 1495 1005 1630
rect 715 1485 755 1495
rect 715 1415 725 1485
rect 745 1415 755 1485
rect 715 1405 755 1415
rect 780 1485 820 1495
rect 780 1415 790 1485
rect 810 1415 820 1485
rect 780 1405 820 1415
rect 845 1485 885 1495
rect 845 1415 855 1485
rect 875 1415 885 1485
rect 845 1405 885 1415
rect 965 1485 1005 1495
rect 965 1415 975 1485
rect 995 1415 1005 1485
rect 965 1405 1005 1415
rect 800 1175 820 1405
rect 965 1380 985 1405
rect 890 1360 985 1380
rect 890 1275 910 1360
rect 930 1330 970 1340
rect 930 1310 940 1330
rect 960 1320 970 1330
rect 960 1310 1010 1320
rect 930 1300 1010 1310
rect 890 1265 970 1275
rect 890 1255 940 1265
rect 930 1245 940 1255
rect 960 1245 970 1265
rect 930 1235 970 1245
rect 990 1215 1010 1300
rect 965 1195 1010 1215
rect 800 1155 880 1175
rect 800 1125 840 1135
rect 800 1115 810 1125
rect 760 1105 810 1115
rect 830 1105 840 1125
rect 760 1095 840 1105
rect 760 1010 780 1095
rect 860 1070 880 1155
rect 800 1060 880 1070
rect 800 1040 810 1060
rect 830 1050 880 1060
rect 830 1040 840 1050
rect 800 1030 840 1040
rect 760 990 800 1010
rect 780 965 800 990
rect 965 965 985 1195
rect 1035 965 1055 1630
rect 1470 1570 1480 1640
rect 1500 1570 1510 1640
rect 1470 1560 1510 1570
rect 1610 1640 1650 1650
rect 1610 1570 1620 1640
rect 1640 1570 1650 1640
rect 1670 1640 1680 1660
rect 1700 1640 1710 1660
rect 1670 1630 1710 1640
rect 1735 1660 1775 1670
rect 1735 1640 1745 1660
rect 1765 1640 1775 1660
rect 2370 1660 2410 1670
rect 1735 1630 1775 1640
rect 2170 1640 2210 1650
rect 1610 1560 1650 1570
rect 1685 1495 1705 1630
rect 1415 1485 1455 1495
rect 1415 1415 1425 1485
rect 1445 1415 1455 1485
rect 1415 1405 1455 1415
rect 1480 1485 1520 1495
rect 1480 1415 1490 1485
rect 1510 1415 1520 1485
rect 1480 1405 1520 1415
rect 1545 1485 1585 1495
rect 1545 1415 1555 1485
rect 1575 1415 1585 1485
rect 1545 1405 1585 1415
rect 1665 1485 1705 1495
rect 1665 1415 1675 1485
rect 1695 1415 1705 1485
rect 1665 1405 1705 1415
rect 1500 1175 1520 1405
rect 1665 1380 1685 1405
rect 1590 1360 1685 1380
rect 1590 1275 1610 1360
rect 1630 1330 1670 1340
rect 1630 1310 1640 1330
rect 1660 1320 1670 1330
rect 1660 1310 1710 1320
rect 1630 1300 1710 1310
rect 1590 1265 1670 1275
rect 1590 1255 1640 1265
rect 1630 1245 1640 1255
rect 1660 1245 1670 1265
rect 1630 1235 1670 1245
rect 1690 1215 1710 1300
rect 1665 1195 1710 1215
rect 1500 1155 1580 1175
rect 1500 1125 1540 1135
rect 1500 1115 1510 1125
rect 1460 1105 1510 1115
rect 1530 1105 1540 1125
rect 1460 1095 1540 1105
rect 1460 1010 1480 1095
rect 1560 1070 1580 1155
rect 1500 1060 1580 1070
rect 1500 1040 1510 1060
rect 1530 1050 1580 1060
rect 1530 1040 1540 1050
rect 1500 1030 1540 1040
rect 1460 990 1500 1010
rect 1480 965 1500 990
rect 1665 965 1685 1195
rect 1735 965 1755 1630
rect 2170 1570 2180 1640
rect 2200 1570 2210 1640
rect 2170 1560 2210 1570
rect 2310 1640 2350 1650
rect 2310 1570 2320 1640
rect 2340 1570 2350 1640
rect 2370 1640 2380 1660
rect 2400 1640 2410 1660
rect 2370 1630 2410 1640
rect 2435 1660 2475 1670
rect 2435 1640 2445 1660
rect 2465 1640 2475 1660
rect 3070 1660 3110 1670
rect 2435 1630 2475 1640
rect 2870 1640 2910 1650
rect 2310 1560 2350 1570
rect 2385 1495 2405 1630
rect 2115 1485 2155 1495
rect 2115 1415 2125 1485
rect 2145 1415 2155 1485
rect 2115 1405 2155 1415
rect 2180 1485 2220 1495
rect 2180 1415 2190 1485
rect 2210 1415 2220 1485
rect 2180 1405 2220 1415
rect 2245 1485 2285 1495
rect 2245 1415 2255 1485
rect 2275 1415 2285 1485
rect 2245 1405 2285 1415
rect 2365 1485 2405 1495
rect 2365 1415 2375 1485
rect 2395 1415 2405 1485
rect 2365 1405 2405 1415
rect 2200 1175 2220 1405
rect 2365 1380 2385 1405
rect 2290 1360 2385 1380
rect 2290 1275 2310 1360
rect 2330 1330 2370 1340
rect 2330 1310 2340 1330
rect 2360 1320 2370 1330
rect 2360 1310 2410 1320
rect 2330 1300 2410 1310
rect 2290 1265 2370 1275
rect 2290 1255 2340 1265
rect 2330 1245 2340 1255
rect 2360 1245 2370 1265
rect 2330 1235 2370 1245
rect 2390 1215 2410 1300
rect 2365 1195 2410 1215
rect 2200 1155 2280 1175
rect 2200 1125 2240 1135
rect 2200 1115 2210 1125
rect 2160 1105 2210 1115
rect 2230 1105 2240 1125
rect 2160 1095 2240 1105
rect 2160 1010 2180 1095
rect 2260 1070 2280 1155
rect 2200 1060 2280 1070
rect 2200 1040 2210 1060
rect 2230 1050 2280 1060
rect 2230 1040 2240 1050
rect 2200 1030 2240 1040
rect 2160 990 2200 1010
rect 2180 965 2200 990
rect 2365 965 2385 1195
rect 2435 965 2455 1630
rect 2870 1570 2880 1640
rect 2900 1570 2910 1640
rect 2870 1560 2910 1570
rect 3010 1640 3050 1650
rect 3010 1570 3020 1640
rect 3040 1570 3050 1640
rect 3070 1640 3080 1660
rect 3100 1640 3110 1660
rect 3070 1630 3110 1640
rect 3135 1660 3175 1670
rect 3135 1640 3145 1660
rect 3165 1640 3175 1660
rect 3770 1660 3810 1670
rect 3135 1630 3175 1640
rect 3570 1640 3610 1650
rect 3010 1560 3050 1570
rect 3085 1495 3105 1630
rect 2815 1485 2855 1495
rect 2815 1415 2825 1485
rect 2845 1415 2855 1485
rect 2815 1405 2855 1415
rect 2880 1485 2920 1495
rect 2880 1415 2890 1485
rect 2910 1415 2920 1485
rect 2880 1405 2920 1415
rect 2945 1485 2985 1495
rect 2945 1415 2955 1485
rect 2975 1415 2985 1485
rect 2945 1405 2985 1415
rect 3065 1485 3105 1495
rect 3065 1415 3075 1485
rect 3095 1415 3105 1485
rect 3065 1405 3105 1415
rect 2900 1175 2920 1405
rect 3065 1380 3085 1405
rect 2990 1360 3085 1380
rect 2990 1275 3010 1360
rect 3030 1330 3070 1340
rect 3030 1310 3040 1330
rect 3060 1320 3070 1330
rect 3060 1310 3110 1320
rect 3030 1300 3110 1310
rect 2990 1265 3070 1275
rect 2990 1255 3040 1265
rect 3030 1245 3040 1255
rect 3060 1245 3070 1265
rect 3030 1235 3070 1245
rect 3090 1215 3110 1300
rect 3065 1195 3110 1215
rect 2900 1155 2980 1175
rect 2900 1125 2940 1135
rect 2900 1115 2910 1125
rect 2860 1105 2910 1115
rect 2930 1105 2940 1125
rect 2860 1095 2940 1105
rect 2860 1010 2880 1095
rect 2960 1070 2980 1155
rect 2900 1060 2980 1070
rect 2900 1040 2910 1060
rect 2930 1050 2980 1060
rect 2930 1040 2940 1050
rect 2900 1030 2940 1040
rect 2860 990 2900 1010
rect 2880 965 2900 990
rect 3065 965 3085 1195
rect 3135 965 3155 1630
rect 3570 1570 3580 1640
rect 3600 1570 3610 1640
rect 3570 1560 3610 1570
rect 3710 1640 3750 1650
rect 3710 1570 3720 1640
rect 3740 1570 3750 1640
rect 3770 1640 3780 1660
rect 3800 1640 3810 1660
rect 3770 1630 3810 1640
rect 3835 1660 3875 1670
rect 3835 1640 3845 1660
rect 3865 1640 3875 1660
rect 4470 1660 4510 1670
rect 3835 1630 3875 1640
rect 4270 1640 4310 1650
rect 3710 1560 3750 1570
rect 3785 1495 3805 1630
rect 3515 1485 3555 1495
rect 3515 1415 3525 1485
rect 3545 1415 3555 1485
rect 3515 1405 3555 1415
rect 3580 1485 3620 1495
rect 3580 1415 3590 1485
rect 3610 1415 3620 1485
rect 3580 1405 3620 1415
rect 3645 1485 3685 1495
rect 3645 1415 3655 1485
rect 3675 1415 3685 1485
rect 3645 1405 3685 1415
rect 3765 1485 3805 1495
rect 3765 1415 3775 1485
rect 3795 1415 3805 1485
rect 3765 1405 3805 1415
rect 3600 1175 3620 1405
rect 3765 1380 3785 1405
rect 3690 1360 3785 1380
rect 3690 1275 3710 1360
rect 3730 1330 3770 1340
rect 3730 1310 3740 1330
rect 3760 1320 3770 1330
rect 3760 1310 3810 1320
rect 3730 1300 3810 1310
rect 3690 1265 3770 1275
rect 3690 1255 3740 1265
rect 3730 1245 3740 1255
rect 3760 1245 3770 1265
rect 3730 1235 3770 1245
rect 3790 1215 3810 1300
rect 3765 1195 3810 1215
rect 3600 1155 3680 1175
rect 3600 1125 3640 1135
rect 3600 1115 3610 1125
rect 3560 1105 3610 1115
rect 3630 1105 3640 1125
rect 3560 1095 3640 1105
rect 3560 1010 3580 1095
rect 3660 1070 3680 1155
rect 3600 1060 3680 1070
rect 3600 1040 3610 1060
rect 3630 1050 3680 1060
rect 3630 1040 3640 1050
rect 3600 1030 3640 1040
rect 3560 990 3600 1010
rect 3580 965 3600 990
rect 3765 965 3785 1195
rect 3835 965 3855 1630
rect 4270 1570 4280 1640
rect 4300 1570 4310 1640
rect 4270 1560 4310 1570
rect 4410 1640 4450 1650
rect 4410 1570 4420 1640
rect 4440 1570 4450 1640
rect 4470 1640 4480 1660
rect 4500 1640 4510 1660
rect 4470 1630 4510 1640
rect 4535 1660 4575 1670
rect 4535 1640 4545 1660
rect 4565 1640 4575 1660
rect 4535 1630 4575 1640
rect 4410 1560 4450 1570
rect 4485 1495 4505 1630
rect 4215 1485 4255 1495
rect 4215 1415 4225 1485
rect 4245 1415 4255 1485
rect 4215 1405 4255 1415
rect 4280 1485 4320 1495
rect 4280 1415 4290 1485
rect 4310 1415 4320 1485
rect 4280 1405 4320 1415
rect 4345 1485 4385 1495
rect 4345 1415 4355 1485
rect 4375 1415 4385 1485
rect 4345 1405 4385 1415
rect 4465 1485 4505 1495
rect 4465 1415 4475 1485
rect 4495 1415 4505 1485
rect 4465 1405 4505 1415
rect 4300 1175 4320 1405
rect 4465 1380 4485 1405
rect 4390 1360 4485 1380
rect 4390 1275 4410 1360
rect 4430 1330 4470 1340
rect 4430 1310 4440 1330
rect 4460 1320 4470 1330
rect 4460 1310 4510 1320
rect 4430 1300 4510 1310
rect 4390 1265 4470 1275
rect 4390 1255 4440 1265
rect 4430 1245 4440 1255
rect 4460 1245 4470 1265
rect 4430 1235 4470 1245
rect 4490 1215 4510 1300
rect 4465 1195 4510 1215
rect 4300 1155 4380 1175
rect 4300 1125 4340 1135
rect 4300 1115 4310 1125
rect 4260 1105 4310 1115
rect 4330 1105 4340 1125
rect 4260 1095 4340 1105
rect 4260 1010 4280 1095
rect 4360 1070 4380 1155
rect 4300 1060 4380 1070
rect 4300 1040 4310 1060
rect 4330 1050 4380 1060
rect 4330 1040 4340 1050
rect 4300 1030 4340 1040
rect 4260 990 4300 1010
rect 4280 965 4300 990
rect 4465 965 4485 1195
rect 4535 965 4555 1630
rect 305 945 355 965
rect 715 955 755 965
rect 715 885 725 955
rect 745 885 755 955
rect 715 875 755 885
rect 780 955 820 965
rect 780 885 790 955
rect 810 885 820 955
rect 780 875 820 885
rect 845 955 885 965
rect 845 885 855 955
rect 875 885 885 955
rect 845 875 885 885
rect 965 955 1055 965
rect 965 885 975 955
rect 995 945 1055 955
rect 1415 955 1455 965
rect 995 885 1005 945
rect 965 875 1005 885
rect 1415 885 1425 955
rect 1445 885 1455 955
rect 1415 875 1455 885
rect 1480 955 1520 965
rect 1480 885 1490 955
rect 1510 885 1520 955
rect 1480 875 1520 885
rect 1545 955 1585 965
rect 1545 885 1555 955
rect 1575 885 1585 955
rect 1545 875 1585 885
rect 1665 955 1755 965
rect 1665 885 1675 955
rect 1695 945 1755 955
rect 2115 955 2155 965
rect 1695 885 1705 945
rect 1665 875 1705 885
rect 2115 885 2125 955
rect 2145 885 2155 955
rect 2115 875 2155 885
rect 2180 955 2220 965
rect 2180 885 2190 955
rect 2210 885 2220 955
rect 2180 875 2220 885
rect 2245 955 2285 965
rect 2245 885 2255 955
rect 2275 885 2285 955
rect 2245 875 2285 885
rect 2365 955 2455 965
rect 2365 885 2375 955
rect 2395 945 2455 955
rect 2815 955 2855 965
rect 2395 885 2405 945
rect 2365 875 2405 885
rect 2815 885 2825 955
rect 2845 885 2855 955
rect 2815 875 2855 885
rect 2880 955 2920 965
rect 2880 885 2890 955
rect 2910 885 2920 955
rect 2880 875 2920 885
rect 2945 955 2985 965
rect 2945 885 2955 955
rect 2975 885 2985 955
rect 2945 875 2985 885
rect 3065 955 3155 965
rect 3065 885 3075 955
rect 3095 945 3155 955
rect 3515 955 3555 965
rect 3095 885 3105 945
rect 3065 875 3105 885
rect 3515 885 3525 955
rect 3545 885 3555 955
rect 3515 875 3555 885
rect 3580 955 3620 965
rect 3580 885 3590 955
rect 3610 885 3620 955
rect 3580 875 3620 885
rect 3645 955 3685 965
rect 3645 885 3655 955
rect 3675 885 3685 955
rect 3645 875 3685 885
rect 3765 955 3855 965
rect 3765 885 3775 955
rect 3795 945 3855 955
rect 4215 955 4255 965
rect 3795 885 3805 945
rect 3765 875 3805 885
rect 4215 885 4225 955
rect 4245 885 4255 955
rect 4215 875 4255 885
rect 4280 955 4320 965
rect 4280 885 4290 955
rect 4310 885 4320 955
rect 4280 875 4320 885
rect 4345 955 4385 965
rect 4345 885 4355 955
rect 4375 885 4385 955
rect 4345 875 4385 885
rect 4465 955 4555 965
rect 4465 885 4475 955
rect 4495 945 4555 955
rect 4495 885 4505 945
rect 4465 875 4505 885
rect 800 815 820 875
rect 965 850 985 875
rect 920 830 985 850
rect 800 795 860 815
rect 840 770 860 795
rect 920 770 940 830
rect 1500 815 1520 875
rect 1665 850 1685 875
rect 1620 830 1685 850
rect 1500 795 1560 815
rect 1540 770 1560 795
rect 1620 770 1640 830
rect 2200 815 2220 875
rect 2365 850 2385 875
rect 2320 830 2385 850
rect 2200 795 2260 815
rect 2240 770 2260 795
rect 2320 770 2340 830
rect 2900 815 2920 875
rect 3065 850 3085 875
rect 3020 830 3085 850
rect 2900 795 2960 815
rect 2940 770 2960 795
rect 3020 770 3040 830
rect 3600 815 3620 875
rect 3765 850 3785 875
rect 3720 830 3785 850
rect 3600 795 3660 815
rect 3640 770 3660 795
rect 3720 770 3740 830
rect 4300 815 4320 875
rect 4465 850 4485 875
rect 4420 830 4485 850
rect 4300 795 4360 815
rect 4340 770 4360 795
rect 4420 770 4440 830
rect 715 760 755 770
rect 715 690 725 760
rect 745 690 755 760
rect 715 680 755 690
rect 820 760 860 770
rect 820 690 830 760
rect 850 690 860 760
rect 820 680 860 690
rect 840 660 860 680
rect 900 760 940 770
rect 900 690 910 760
rect 930 690 940 760
rect 900 680 940 690
rect 965 760 1005 770
rect 965 690 975 760
rect 995 690 1005 760
rect 965 680 1005 690
rect 1415 760 1455 770
rect 1415 690 1425 760
rect 1445 690 1455 760
rect 1415 680 1455 690
rect 1520 760 1560 770
rect 1520 690 1530 760
rect 1550 690 1560 760
rect 1520 680 1560 690
rect 840 640 880 660
rect 800 610 840 620
rect 800 600 810 610
rect 760 590 810 600
rect 830 590 840 610
rect 760 580 840 590
rect 760 495 780 580
rect 860 555 880 640
rect 800 545 880 555
rect 800 525 810 545
rect 830 535 880 545
rect 830 525 840 535
rect 800 515 840 525
rect 760 475 840 495
rect 820 280 840 475
rect 900 405 920 680
rect 1540 660 1560 680
rect 1600 760 1640 770
rect 1600 690 1610 760
rect 1630 690 1640 760
rect 1600 680 1640 690
rect 1665 760 1705 770
rect 1665 690 1675 760
rect 1695 690 1705 760
rect 1665 680 1705 690
rect 2115 760 2155 770
rect 2115 690 2125 760
rect 2145 690 2155 760
rect 2115 680 2155 690
rect 2220 760 2260 770
rect 2220 690 2230 760
rect 2250 690 2260 760
rect 2220 680 2260 690
rect 1540 640 1580 660
rect 1500 610 1540 620
rect 1500 600 1510 610
rect 1460 590 1510 600
rect 1530 590 1540 610
rect 1460 580 1540 590
rect 1460 495 1480 580
rect 1560 555 1580 640
rect 1500 545 1580 555
rect 1500 525 1510 545
rect 1530 535 1580 545
rect 1530 525 1540 535
rect 1500 515 1540 525
rect 1460 475 1540 495
rect 940 455 980 465
rect 940 435 950 455
rect 970 445 980 455
rect 970 435 1000 445
rect 940 425 1000 435
rect 900 385 940 405
rect 920 375 960 385
rect 920 355 930 375
rect 950 355 960 375
rect 920 345 960 355
rect 980 320 1000 425
rect 920 300 1000 320
rect 920 280 940 300
rect 1520 280 1540 475
rect 1600 405 1620 680
rect 2240 660 2260 680
rect 2300 760 2340 770
rect 2300 690 2310 760
rect 2330 690 2340 760
rect 2300 680 2340 690
rect 2365 760 2405 770
rect 2365 690 2375 760
rect 2395 690 2405 760
rect 2365 680 2405 690
rect 2815 760 2855 770
rect 2815 690 2825 760
rect 2845 690 2855 760
rect 2815 680 2855 690
rect 2920 760 2960 770
rect 2920 690 2930 760
rect 2950 690 2960 760
rect 2920 680 2960 690
rect 2240 640 2280 660
rect 2200 610 2240 620
rect 2200 600 2210 610
rect 2160 590 2210 600
rect 2230 590 2240 610
rect 2160 580 2240 590
rect 2160 495 2180 580
rect 2260 555 2280 640
rect 2200 545 2280 555
rect 2200 525 2210 545
rect 2230 535 2280 545
rect 2230 525 2240 535
rect 2200 515 2240 525
rect 2160 475 2240 495
rect 1640 455 1680 465
rect 1640 435 1650 455
rect 1670 445 1680 455
rect 1670 435 1700 445
rect 1640 425 1700 435
rect 1600 385 1640 405
rect 1620 375 1660 385
rect 1620 355 1630 375
rect 1650 355 1660 375
rect 1620 345 1660 355
rect 1680 320 1700 425
rect 1620 300 1700 320
rect 1620 280 1640 300
rect 2220 280 2240 475
rect 2300 405 2320 680
rect 2940 660 2960 680
rect 3000 760 3040 770
rect 3000 690 3010 760
rect 3030 690 3040 760
rect 3000 680 3040 690
rect 3065 760 3105 770
rect 3065 690 3075 760
rect 3095 690 3105 760
rect 3065 680 3105 690
rect 3515 760 3555 770
rect 3515 690 3525 760
rect 3545 690 3555 760
rect 3515 680 3555 690
rect 3620 760 3660 770
rect 3620 690 3630 760
rect 3650 690 3660 760
rect 3620 680 3660 690
rect 2940 640 2980 660
rect 2900 610 2940 620
rect 2900 600 2910 610
rect 2860 590 2910 600
rect 2930 590 2940 610
rect 2860 580 2940 590
rect 2860 495 2880 580
rect 2960 555 2980 640
rect 2900 545 2980 555
rect 2900 525 2910 545
rect 2930 535 2980 545
rect 2930 525 2940 535
rect 2900 515 2940 525
rect 2860 475 2940 495
rect 2340 455 2380 465
rect 2340 435 2350 455
rect 2370 445 2380 455
rect 2370 435 2400 445
rect 2340 425 2400 435
rect 2300 385 2340 405
rect 2320 375 2360 385
rect 2320 355 2330 375
rect 2350 355 2360 375
rect 2320 345 2360 355
rect 2380 320 2400 425
rect 2320 300 2400 320
rect 2320 280 2340 300
rect 2920 280 2940 475
rect 3000 405 3020 680
rect 3640 660 3660 680
rect 3700 760 3740 770
rect 3700 690 3710 760
rect 3730 690 3740 760
rect 3700 680 3740 690
rect 3765 760 3805 770
rect 3765 690 3775 760
rect 3795 690 3805 760
rect 3765 680 3805 690
rect 4215 760 4255 770
rect 4215 690 4225 760
rect 4245 690 4255 760
rect 4215 680 4255 690
rect 4320 760 4360 770
rect 4320 690 4330 760
rect 4350 690 4360 760
rect 4320 680 4360 690
rect 3640 640 3680 660
rect 3600 610 3640 620
rect 3600 600 3610 610
rect 3560 590 3610 600
rect 3630 590 3640 610
rect 3560 580 3640 590
rect 3560 495 3580 580
rect 3660 555 3680 640
rect 3600 545 3680 555
rect 3600 525 3610 545
rect 3630 535 3680 545
rect 3630 525 3640 535
rect 3600 515 3640 525
rect 3560 475 3640 495
rect 3040 455 3080 465
rect 3040 435 3050 455
rect 3070 445 3080 455
rect 3070 435 3100 445
rect 3040 425 3100 435
rect 3000 385 3040 405
rect 3020 375 3060 385
rect 3020 355 3030 375
rect 3050 355 3060 375
rect 3020 345 3060 355
rect 3080 320 3100 425
rect 3020 300 3100 320
rect 3020 280 3040 300
rect 3620 280 3640 475
rect 3700 405 3720 680
rect 4340 660 4360 680
rect 4400 760 4440 770
rect 4400 690 4410 760
rect 4430 690 4440 760
rect 4400 680 4440 690
rect 4465 760 4505 770
rect 4465 690 4475 760
rect 4495 690 4505 760
rect 4465 680 4505 690
rect 4340 640 4380 660
rect 4300 610 4340 620
rect 4300 600 4310 610
rect 4260 590 4310 600
rect 4330 590 4340 610
rect 4260 580 4340 590
rect 4260 495 4280 580
rect 4360 555 4380 640
rect 4300 545 4380 555
rect 4300 525 4310 545
rect 4330 535 4380 545
rect 4330 525 4340 535
rect 4300 515 4340 525
rect 4260 475 4340 495
rect 3740 455 3780 465
rect 3740 435 3750 455
rect 3770 445 3780 455
rect 3770 435 3800 445
rect 3740 425 3800 435
rect 3700 385 3740 405
rect 3720 375 3760 385
rect 3720 355 3730 375
rect 3750 355 3760 375
rect 3720 345 3760 355
rect 3780 320 3800 425
rect 3720 300 3800 320
rect 3720 280 3740 300
rect 4320 280 4340 475
rect 4400 405 4420 680
rect 4440 455 4480 465
rect 4440 435 4450 455
rect 4470 445 4480 455
rect 4470 435 4500 445
rect 4440 425 4500 435
rect 4400 385 4440 405
rect 4420 375 4460 385
rect 4420 355 4430 375
rect 4450 355 4460 375
rect 4420 345 4460 355
rect 4480 320 4500 425
rect 4420 300 4500 320
rect 4420 280 4440 300
rect 715 270 755 280
rect 715 200 725 270
rect 745 200 755 270
rect 715 190 755 200
rect 820 270 860 280
rect 820 200 830 270
rect 850 200 860 270
rect 820 190 860 200
rect 900 270 940 280
rect 900 200 910 270
rect 930 200 940 270
rect 900 190 940 200
rect 965 270 1005 280
rect 965 200 975 270
rect 995 200 1005 270
rect 965 190 1005 200
rect 1415 270 1455 280
rect 1415 200 1425 270
rect 1445 200 1455 270
rect 1415 190 1455 200
rect 1520 270 1560 280
rect 1520 200 1530 270
rect 1550 200 1560 270
rect 1520 190 1560 200
rect 1600 270 1640 280
rect 1600 200 1610 270
rect 1630 200 1640 270
rect 1600 190 1640 200
rect 1665 270 1705 280
rect 1665 200 1675 270
rect 1695 200 1705 270
rect 1665 190 1705 200
rect 2115 270 2155 280
rect 2115 200 2125 270
rect 2145 200 2155 270
rect 2115 190 2155 200
rect 2220 270 2260 280
rect 2220 200 2230 270
rect 2250 200 2260 270
rect 2220 190 2260 200
rect 2300 270 2340 280
rect 2300 200 2310 270
rect 2330 200 2340 270
rect 2300 190 2340 200
rect 2365 270 2405 280
rect 2365 200 2375 270
rect 2395 200 2405 270
rect 2365 190 2405 200
rect 2815 270 2855 280
rect 2815 200 2825 270
rect 2845 200 2855 270
rect 2815 190 2855 200
rect 2920 270 2960 280
rect 2920 200 2930 270
rect 2950 200 2960 270
rect 2920 190 2960 200
rect 3000 270 3040 280
rect 3000 200 3010 270
rect 3030 200 3040 270
rect 3000 190 3040 200
rect 3065 270 3105 280
rect 3065 200 3075 270
rect 3095 200 3105 270
rect 3065 190 3105 200
rect 3515 270 3555 280
rect 3515 200 3525 270
rect 3545 200 3555 270
rect 3515 190 3555 200
rect 3620 270 3660 280
rect 3620 200 3630 270
rect 3650 200 3660 270
rect 3620 190 3660 200
rect 3700 270 3740 280
rect 3700 200 3710 270
rect 3730 200 3740 270
rect 3700 190 3740 200
rect 3765 270 3805 280
rect 3765 200 3775 270
rect 3795 200 3805 270
rect 3765 190 3805 200
rect 4215 270 4255 280
rect 4215 200 4225 270
rect 4245 200 4255 270
rect 4215 190 4255 200
rect 4320 270 4360 280
rect 4320 200 4330 270
rect 4350 200 4360 270
rect 4320 190 4360 200
rect 4400 270 4440 280
rect 4400 200 4410 270
rect 4430 200 4440 270
rect 4400 190 4440 200
rect 4465 270 4505 280
rect 4465 200 4475 270
rect 4495 200 4505 270
rect 4465 190 4505 200
rect 790 140 830 150
rect 790 70 800 140
rect 820 70 830 140
rect 790 60 830 70
rect 925 140 965 150
rect 925 70 935 140
rect 955 70 965 140
rect 925 60 965 70
rect 1490 140 1530 150
rect 1490 70 1500 140
rect 1520 70 1530 140
rect 1490 60 1530 70
rect 1625 140 1665 150
rect 1625 70 1635 140
rect 1655 70 1665 140
rect 1625 60 1665 70
rect 2190 140 2230 150
rect 2190 70 2200 140
rect 2220 70 2230 140
rect 2190 60 2230 70
rect 2325 140 2365 150
rect 2325 70 2335 140
rect 2355 70 2365 140
rect 2325 60 2365 70
rect 2890 140 2930 150
rect 2890 70 2900 140
rect 2920 70 2930 140
rect 2890 60 2930 70
rect 3025 140 3065 150
rect 3025 70 3035 140
rect 3055 70 3065 140
rect 3025 60 3065 70
rect 3590 140 3630 150
rect 3590 70 3600 140
rect 3620 70 3630 140
rect 3590 60 3630 70
rect 3725 140 3765 150
rect 3725 70 3735 140
rect 3755 70 3765 140
rect 3725 60 3765 70
rect 4290 140 4330 150
rect 4290 70 4300 140
rect 4320 70 4330 140
rect 4290 60 4330 70
rect 4425 140 4465 150
rect 4425 70 4435 140
rect 4455 70 4465 140
rect 4425 60 4465 70
rect 735 30 775 40
rect 735 10 745 30
rect 765 10 775 30
rect 735 0 775 10
rect 855 30 895 40
rect 855 10 865 30
rect 885 10 895 30
rect 855 0 895 10
rect 1435 30 1475 40
rect 1435 10 1445 30
rect 1465 10 1475 30
rect 1435 0 1475 10
rect 1555 30 1595 40
rect 1555 10 1565 30
rect 1585 10 1595 30
rect 1555 0 1595 10
rect 2135 30 2175 40
rect 2135 10 2145 30
rect 2165 10 2175 30
rect 2135 0 2175 10
rect 2255 30 2295 40
rect 2255 10 2265 30
rect 2285 10 2295 30
rect 2255 0 2295 10
rect 2835 30 2875 40
rect 2835 10 2845 30
rect 2865 10 2875 30
rect 2835 0 2875 10
rect 2955 30 2995 40
rect 2955 10 2965 30
rect 2985 10 2995 30
rect 2955 0 2995 10
rect 3535 30 3575 40
rect 3535 10 3545 30
rect 3565 10 3575 30
rect 3535 0 3575 10
rect 3655 30 3695 40
rect 3655 10 3665 30
rect 3685 10 3695 30
rect 3655 0 3695 10
rect 4235 30 4275 40
rect 4235 10 4245 30
rect 4265 10 4275 30
rect 4235 0 4275 10
rect 4355 30 4395 40
rect 4355 10 4365 30
rect 4385 10 4395 30
rect 4355 0 4395 10
<< viali >>
rect 780 1570 800 1640
rect 920 1570 940 1640
rect 855 1415 875 1485
rect 1480 1570 1500 1640
rect 1620 1570 1640 1640
rect 1555 1415 1575 1485
rect 2180 1570 2200 1640
rect 2320 1570 2340 1640
rect 2255 1415 2275 1485
rect 2880 1570 2900 1640
rect 3020 1570 3040 1640
rect 2955 1415 2975 1485
rect 3580 1570 3600 1640
rect 3720 1570 3740 1640
rect 3655 1415 3675 1485
rect 4280 1570 4300 1640
rect 4420 1570 4440 1640
rect 4355 1415 4375 1485
rect 855 885 875 955
rect 1555 885 1575 955
rect 2255 885 2275 955
rect 2955 885 2975 955
rect 3655 885 3675 955
rect 4355 885 4375 955
rect 725 690 745 760
rect 975 690 995 760
rect 1425 690 1445 760
rect 1675 690 1695 760
rect 2125 690 2145 760
rect 2375 690 2395 760
rect 2825 690 2845 760
rect 3075 690 3095 760
rect 3525 690 3545 760
rect 3775 690 3795 760
rect 4225 690 4245 760
rect 4475 690 4495 760
rect 725 200 745 270
rect 975 200 995 270
rect 1425 200 1445 270
rect 1675 200 1695 270
rect 2125 200 2145 270
rect 2375 200 2395 270
rect 2825 200 2845 270
rect 3075 200 3095 270
rect 3525 200 3545 270
rect 3775 200 3795 270
rect 4225 200 4245 270
rect 4475 200 4495 270
rect 800 70 820 140
rect 935 70 955 140
rect 1500 70 1520 140
rect 1635 70 1655 140
rect 2200 70 2220 140
rect 2335 70 2355 140
rect 2900 70 2920 140
rect 3035 70 3055 140
rect 3600 70 3620 140
rect 3735 70 3755 140
rect 4300 70 4320 140
rect 4435 70 4455 140
rect 745 10 765 30
rect 865 10 885 30
rect 1445 10 1465 30
rect 1565 10 1585 30
rect 2145 10 2165 30
rect 2265 10 2285 30
rect 2845 10 2865 30
rect 2965 10 2985 30
rect 3545 10 3565 30
rect 3665 10 3685 30
rect 4245 10 4265 30
rect 4365 10 4385 30
<< metal1 >>
rect 330 1640 4610 1675
rect 330 1570 780 1640
rect 800 1570 920 1640
rect 940 1570 1480 1640
rect 1500 1570 1620 1640
rect 1640 1570 2180 1640
rect 2200 1570 2320 1640
rect 2340 1570 2880 1640
rect 2900 1570 3020 1640
rect 3040 1570 3580 1640
rect 3600 1570 3720 1640
rect 3740 1570 4280 1640
rect 4300 1570 4420 1640
rect 4440 1570 4610 1640
rect 330 1540 4610 1570
rect 330 1535 415 1540
rect 690 1535 4610 1540
rect 845 1485 885 1535
rect 845 1415 855 1485
rect 875 1415 885 1485
rect 845 955 885 1415
rect 845 885 855 955
rect 875 885 885 955
rect 845 875 885 885
rect 1545 1485 1585 1535
rect 1545 1415 1555 1485
rect 1575 1415 1585 1485
rect 1545 955 1585 1415
rect 1545 885 1555 955
rect 1575 885 1585 955
rect 1545 875 1585 885
rect 2245 1485 2285 1535
rect 2245 1415 2255 1485
rect 2275 1415 2285 1485
rect 2245 955 2285 1415
rect 2245 885 2255 955
rect 2275 885 2285 955
rect 2245 875 2285 885
rect 2945 1485 2985 1535
rect 2945 1415 2955 1485
rect 2975 1415 2985 1485
rect 2945 955 2985 1415
rect 2945 885 2955 955
rect 2975 885 2985 955
rect 2945 875 2985 885
rect 3645 1485 3685 1535
rect 3645 1415 3655 1485
rect 3675 1415 3685 1485
rect 3645 955 3685 1415
rect 3645 885 3655 955
rect 3675 885 3685 955
rect 3645 875 3685 885
rect 4345 1485 4385 1535
rect 4345 1415 4355 1485
rect 4375 1415 4385 1485
rect 4345 955 4385 1415
rect 4345 885 4355 955
rect 4375 885 4385 955
rect 4345 875 4385 885
rect 310 760 755 775
rect 310 690 725 760
rect 745 690 755 760
rect 310 675 755 690
rect 710 270 755 675
rect 710 200 725 270
rect 745 200 755 270
rect 710 155 755 200
rect 965 760 1455 775
rect 965 690 975 760
rect 995 690 1425 760
rect 1445 690 1455 760
rect 965 675 1455 690
rect 965 270 1010 675
rect 965 200 975 270
rect 995 200 1010 270
rect 965 155 1010 200
rect 1410 270 1455 675
rect 1410 200 1425 270
rect 1445 200 1455 270
rect 1410 155 1455 200
rect 1665 760 2155 775
rect 1665 690 1675 760
rect 1695 690 2125 760
rect 2145 690 2155 760
rect 1665 675 2155 690
rect 1665 270 1710 675
rect 1665 200 1675 270
rect 1695 200 1710 270
rect 1665 155 1710 200
rect 2110 270 2155 675
rect 2110 200 2125 270
rect 2145 200 2155 270
rect 2110 155 2155 200
rect 2365 760 2855 775
rect 2365 690 2375 760
rect 2395 690 2825 760
rect 2845 690 2855 760
rect 2365 675 2855 690
rect 2365 270 2410 675
rect 2365 200 2375 270
rect 2395 200 2410 270
rect 2365 155 2410 200
rect 2810 270 2855 675
rect 2810 200 2825 270
rect 2845 200 2855 270
rect 2810 155 2855 200
rect 3065 760 3555 775
rect 3065 690 3075 760
rect 3095 690 3525 760
rect 3545 690 3555 760
rect 3065 675 3555 690
rect 3065 270 3110 675
rect 3065 200 3075 270
rect 3095 200 3110 270
rect 3065 155 3110 200
rect 3510 270 3555 675
rect 3510 200 3525 270
rect 3545 200 3555 270
rect 3510 155 3555 200
rect 3765 760 4255 775
rect 3765 690 3775 760
rect 3795 690 4225 760
rect 4245 690 4255 760
rect 3765 675 4255 690
rect 3765 270 3810 675
rect 3765 200 3775 270
rect 3795 200 3810 270
rect 3765 155 3810 200
rect 4210 270 4255 675
rect 4210 200 4225 270
rect 4245 200 4255 270
rect 4210 155 4255 200
rect 4465 760 4535 775
rect 4465 690 4475 760
rect 4495 690 4535 760
rect 4465 675 4535 690
rect 4465 270 4510 675
rect 4465 200 4475 270
rect 4495 200 4510 270
rect 4465 155 4510 200
rect 310 140 4535 155
rect 310 70 800 140
rect 820 70 935 140
rect 955 70 1500 140
rect 1520 70 1635 140
rect 1655 70 2200 140
rect 2220 70 2335 140
rect 2355 70 2900 140
rect 2920 70 3035 140
rect 3055 70 3600 140
rect 3620 70 3735 140
rect 3755 70 4300 140
rect 4320 70 4435 140
rect 4455 70 4535 140
rect 310 55 4535 70
rect 310 30 4535 40
rect 310 10 745 30
rect 765 10 865 30
rect 885 10 1445 30
rect 1465 10 1565 30
rect 1585 10 2145 30
rect 2165 10 2265 30
rect 2285 10 2845 30
rect 2865 10 2965 30
rect 2985 10 3545 30
rect 3565 10 3665 30
rect 3685 10 4245 30
rect 4265 10 4365 30
rect 4385 10 4535 30
rect 310 0 4535 10
use CSRL_latch  CSRL_latch_0 ~/MADVLSI/Miniproject2/layout
timestamp 1699199846
transform 1 0 125 0 1 -490
box -135 490 205 2165
<< labels >>
rlabel metal1 710 20 710 20 7 CLK
port 1 w
rlabel locali 1005 920 1005 920 3 Qn
port 7 e
rlabel pdiff 1010 1450 1010 1450 3 Q
port 6 e
rlabel pdiff 710 920 710 920 7 Dn
port 5 w
rlabel pdiff 710 1450 710 1450 7 D
port 4 w
rlabel metal1 710 105 710 105 7 GND
port 3 w
rlabel metal1 690 1605 690 1605 7 VDD
port 2 w
rlabel poly 1065 1680 1065 1680 5 D0b
port 6 s
rlabel metal1 1410 20 1410 20 7 CLK
port 1 w
rlabel locali 1705 920 1705 920 3 Qn
port 7 e
rlabel pdiff 1710 1450 1710 1450 3 Q
port 6 e
rlabel pdiff 1410 920 1410 920 7 Dn
port 5 w
rlabel pdiff 1410 1450 1410 1450 7 D
port 4 w
rlabel metal1 1410 105 1410 105 7 GND
port 3 w
rlabel metal1 1390 1605 1390 1605 7 VDD
port 2 w
rlabel poly 2465 1680 2465 1680 5 D1b
port 8 s
rlabel poly 2365 1680 2365 1680 5 D1
port 7 s
rlabel poly 1765 1680 1765 1680 5 D0b
port 6 s
rlabel poly 1665 1680 1665 1680 5 D0
port 5 s
rlabel metal1 2110 20 2110 20 7 CLK
port 1 w
rlabel locali 2405 920 2405 920 3 Qn
port 7 e
rlabel pdiff 2410 1450 2410 1450 3 Q
port 6 e
rlabel pdiff 2110 920 2110 920 7 Dn
port 5 w
rlabel pdiff 2110 1450 2110 1450 7 D
port 4 w
rlabel metal1 2110 105 2110 105 7 GND
port 3 w
rlabel metal1 2090 1605 2090 1605 7 VDD
port 2 w
rlabel poly 2465 1680 2465 1680 5 D0b
port 6 s
rlabel poly 2365 1680 2365 1680 5 D0
port 5 s
rlabel metal1 2810 20 2810 20 7 CLK
port 1 w
rlabel locali 3105 920 3105 920 3 Qn
port 7 e
rlabel pdiff 3110 1450 3110 1450 3 Q
port 6 e
rlabel pdiff 2810 920 2810 920 7 Dn
port 5 w
rlabel pdiff 2810 1450 2810 1450 7 D
port 4 w
rlabel metal1 2810 105 2810 105 7 GND
port 3 w
rlabel metal1 2790 1605 2790 1605 7 VDD
port 2 w
rlabel poly 3865 1680 3865 1680 5 D1b
port 8 s
rlabel poly 3765 1680 3765 1680 5 D1
port 7 s
rlabel poly 3165 1680 3165 1680 5 D0b
port 6 s
rlabel poly 3065 1680 3065 1680 5 D0
port 5 s
rlabel metal1 3510 20 3510 20 7 CLK
port 1 w
rlabel locali 3805 920 3805 920 3 Qn
port 7 e
rlabel pdiff 3810 1450 3810 1450 3 Q
port 6 e
rlabel pdiff 3510 920 3510 920 7 Dn
port 5 w
rlabel pdiff 3510 1450 3510 1450 7 D
port 4 w
rlabel metal1 3510 105 3510 105 7 GND
port 3 w
rlabel metal1 3490 1605 3490 1605 7 VDD
port 2 w
rlabel poly 3865 1680 3865 1680 5 D0b
port 6 s
rlabel poly 3765 1680 3765 1680 5 D0
port 5 s
rlabel metal1 4210 20 4210 20 7 CLK
port 1 w
rlabel locali 4505 920 4505 920 3 Qn
port 7 e
rlabel pdiff 4510 1450 4510 1450 3 Q
port 6 e
rlabel pdiff 4210 920 4210 920 7 Dn
port 5 w
rlabel pdiff 4210 1450 4210 1450 7 D
port 4 w
rlabel metal1 4210 105 4210 105 7 GND
port 3 w
rlabel metal1 4190 1605 4190 1605 7 VDD
port 2 w
rlabel poly 4565 1680 4565 1680 5 D0b
port 6 s
rlabel poly 4465 1680 4465 1680 5 D0
port 5 s
<< end >>

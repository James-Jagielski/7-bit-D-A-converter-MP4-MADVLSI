magic
tech sky130A
timestamp 1699140029
<< locali >>
rect 340 1500 360 1680
rect 315 1480 360 1500
rect 315 1410 340 1430
rect 320 1390 340 1410
rect 320 1380 360 1390
rect 320 1360 330 1380
rect 350 1360 360 1380
rect 320 1350 360 1360
rect 380 970 400 1680
rect 420 1380 460 1390
rect 420 1360 430 1380
rect 450 1360 460 1380
rect 420 1350 460 1360
rect 315 950 425 970
rect 315 685 425 715
rect 315 195 425 225
<< viali >>
rect 330 1360 350 1380
rect 430 1360 450 1380
<< metal1 >>
rect 340 1540 425 1680
rect 320 1380 460 1390
rect 320 1360 330 1380
rect 350 1360 430 1380
rect 450 1360 460 1380
rect 320 1350 460 1360
rect 320 60 425 160
rect 320 5 425 45
use CSRL_latch  CSRL_latch_0 ~/MADVLSI/Miniproject2/layout
timestamp 1699138609
transform 1 0 135 0 1 -485
box -135 490 205 2165
<< end >>

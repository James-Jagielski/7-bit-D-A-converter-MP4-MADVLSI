magic
tech sky130A
timestamp 1699928585
<< nwell >>
rect -110 690 1880 1400
<< nmos >>
rect 10 10 60 610
rect 110 10 160 610
rect 210 10 260 610
rect 310 10 360 610
rect 410 10 460 610
rect 610 10 660 610
rect 710 10 760 610
rect 810 10 860 610
rect 910 10 960 610
rect 1110 10 1160 610
rect 1210 10 1260 610
rect 1310 10 1360 610
rect 1410 10 1460 610
rect 1510 10 1560 610
<< pmos >>
rect 10 745 60 1345
rect 110 745 160 1345
rect 210 745 260 1345
rect 310 745 360 1345
rect 410 745 460 1345
rect 610 745 660 1345
rect 710 745 760 1345
rect 810 745 860 1345
rect 910 745 960 1345
rect 1010 745 1060 1345
rect 1110 745 1160 1345
rect 1310 745 1360 1345
rect 1410 745 1460 1345
rect 1510 745 1560 1345
rect 1610 745 1660 1345
rect 1710 745 1760 1345
<< ndiff >>
rect -40 595 10 610
rect -40 320 -25 595
rect -5 320 10 595
rect -40 300 10 320
rect -40 25 -25 300
rect -5 25 10 300
rect -40 10 10 25
rect 60 595 110 610
rect 60 320 75 595
rect 95 320 110 595
rect 60 300 110 320
rect 60 25 75 300
rect 95 25 110 300
rect 60 10 110 25
rect 160 595 210 610
rect 160 320 175 595
rect 195 320 210 595
rect 160 300 210 320
rect 160 25 175 300
rect 195 25 210 300
rect 160 10 210 25
rect 260 595 310 610
rect 260 320 275 595
rect 295 320 310 595
rect 260 300 310 320
rect 260 25 275 300
rect 295 25 310 300
rect 260 10 310 25
rect 360 595 410 610
rect 360 320 375 595
rect 395 320 410 595
rect 360 300 410 320
rect 360 25 375 300
rect 395 25 410 300
rect 360 10 410 25
rect 460 595 510 610
rect 560 595 610 610
rect 460 320 475 595
rect 495 320 510 595
rect 560 320 575 595
rect 595 320 610 595
rect 460 300 510 320
rect 560 300 610 320
rect 460 25 475 300
rect 495 25 510 300
rect 560 25 575 300
rect 595 25 610 300
rect 460 10 510 25
rect 560 10 610 25
rect 660 595 710 610
rect 660 320 675 595
rect 695 320 710 595
rect 660 300 710 320
rect 660 25 675 300
rect 695 25 710 300
rect 660 10 710 25
rect 760 595 810 610
rect 760 320 775 595
rect 795 320 810 595
rect 760 300 810 320
rect 760 25 775 300
rect 795 25 810 300
rect 760 10 810 25
rect 860 595 910 610
rect 860 320 875 595
rect 895 320 910 595
rect 860 300 910 320
rect 860 25 875 300
rect 895 25 910 300
rect 860 10 910 25
rect 960 595 1010 610
rect 1060 595 1110 610
rect 960 320 975 595
rect 995 320 1010 595
rect 1060 320 1075 595
rect 1095 320 1110 595
rect 960 300 1010 320
rect 1060 300 1110 320
rect 960 25 975 300
rect 995 25 1010 300
rect 1060 25 1075 300
rect 1095 25 1110 300
rect 960 10 1010 25
rect 1060 10 1110 25
rect 1160 595 1210 610
rect 1160 320 1175 595
rect 1195 320 1210 595
rect 1160 300 1210 320
rect 1160 25 1175 300
rect 1195 25 1210 300
rect 1160 10 1210 25
rect 1260 595 1310 610
rect 1260 320 1275 595
rect 1295 320 1310 595
rect 1260 300 1310 320
rect 1260 25 1275 300
rect 1295 25 1310 300
rect 1260 10 1310 25
rect 1360 595 1410 610
rect 1360 320 1375 595
rect 1395 320 1410 595
rect 1360 300 1410 320
rect 1360 25 1375 300
rect 1395 25 1410 300
rect 1360 10 1410 25
rect 1460 595 1510 610
rect 1460 320 1475 595
rect 1495 320 1510 595
rect 1460 300 1510 320
rect 1460 25 1475 300
rect 1495 25 1510 300
rect 1460 10 1510 25
rect 1560 595 1610 610
rect 1560 320 1575 595
rect 1595 320 1610 595
rect 1560 300 1610 320
rect 1560 25 1575 300
rect 1595 25 1610 300
rect 1560 10 1610 25
<< pdiff >>
rect -40 1330 10 1345
rect -40 1055 -25 1330
rect -5 1055 10 1330
rect -40 1035 10 1055
rect -40 760 -25 1035
rect -5 760 10 1035
rect -40 745 10 760
rect 60 1330 110 1345
rect 60 1055 75 1330
rect 95 1055 110 1330
rect 60 1035 110 1055
rect 60 760 75 1035
rect 95 760 110 1035
rect 60 745 110 760
rect 160 1330 210 1345
rect 160 1055 175 1330
rect 195 1055 210 1330
rect 160 1035 210 1055
rect 160 760 175 1035
rect 195 760 210 1035
rect 160 745 210 760
rect 260 1330 310 1345
rect 260 1055 275 1330
rect 295 1055 310 1330
rect 260 1035 310 1055
rect 260 760 275 1035
rect 295 760 310 1035
rect 260 745 310 760
rect 360 1330 410 1345
rect 360 1055 375 1330
rect 395 1055 410 1330
rect 360 1035 410 1055
rect 360 760 375 1035
rect 395 760 410 1035
rect 360 745 410 760
rect 460 1330 510 1345
rect 560 1330 610 1345
rect 460 1055 475 1330
rect 495 1055 510 1330
rect 560 1055 575 1330
rect 595 1055 610 1330
rect 460 1035 510 1055
rect 560 1035 610 1055
rect 460 760 475 1035
rect 495 760 510 1035
rect 560 760 575 1035
rect 595 760 610 1035
rect 460 745 510 760
rect 560 745 610 760
rect 660 1330 710 1345
rect 660 1055 675 1330
rect 695 1055 710 1330
rect 660 1035 710 1055
rect 660 760 675 1035
rect 695 760 710 1035
rect 660 745 710 760
rect 760 1330 810 1345
rect 760 1055 775 1330
rect 795 1055 810 1330
rect 760 1035 810 1055
rect 760 760 775 1035
rect 795 760 810 1035
rect 760 745 810 760
rect 860 1330 910 1345
rect 860 1055 875 1330
rect 895 1055 910 1330
rect 860 1035 910 1055
rect 860 760 875 1035
rect 895 760 910 1035
rect 860 745 910 760
rect 960 1330 1010 1345
rect 960 1055 975 1330
rect 995 1055 1010 1330
rect 960 1035 1010 1055
rect 960 760 975 1035
rect 995 760 1010 1035
rect 960 745 1010 760
rect 1060 1330 1110 1345
rect 1060 1055 1075 1330
rect 1095 1055 1110 1330
rect 1060 1035 1110 1055
rect 1060 760 1075 1035
rect 1095 760 1110 1035
rect 1060 745 1110 760
rect 1160 1330 1210 1345
rect 1260 1330 1310 1345
rect 1160 1055 1175 1330
rect 1195 1055 1210 1330
rect 1260 1055 1275 1330
rect 1295 1055 1310 1330
rect 1160 1035 1210 1055
rect 1260 1035 1310 1055
rect 1160 760 1175 1035
rect 1195 760 1210 1035
rect 1260 760 1275 1035
rect 1295 760 1310 1035
rect 1160 745 1210 760
rect 1260 745 1310 760
rect 1360 1330 1410 1345
rect 1360 1055 1375 1330
rect 1395 1055 1410 1330
rect 1360 1035 1410 1055
rect 1360 760 1375 1035
rect 1395 760 1410 1035
rect 1360 745 1410 760
rect 1460 1330 1510 1345
rect 1460 1055 1475 1330
rect 1495 1055 1510 1330
rect 1460 1035 1510 1055
rect 1460 760 1475 1035
rect 1495 760 1510 1035
rect 1460 745 1510 760
rect 1560 1330 1610 1345
rect 1560 1055 1575 1330
rect 1595 1055 1610 1330
rect 1560 1035 1610 1055
rect 1560 760 1575 1035
rect 1595 760 1610 1035
rect 1560 745 1610 760
rect 1660 1330 1710 1345
rect 1660 1055 1675 1330
rect 1695 1055 1710 1330
rect 1660 1035 1710 1055
rect 1660 760 1675 1035
rect 1695 760 1710 1035
rect 1660 745 1710 760
rect 1760 1330 1810 1345
rect 1760 1055 1775 1330
rect 1795 1055 1810 1330
rect 1760 1035 1810 1055
rect 1760 760 1775 1035
rect 1795 760 1810 1035
rect 1760 745 1810 760
<< ndiffc >>
rect -25 320 -5 595
rect -25 25 -5 300
rect 75 320 95 595
rect 75 25 95 300
rect 175 320 195 595
rect 175 25 195 300
rect 275 320 295 595
rect 275 25 295 300
rect 375 320 395 595
rect 375 25 395 300
rect 475 320 495 595
rect 575 320 595 595
rect 475 25 495 300
rect 575 25 595 300
rect 675 320 695 595
rect 675 25 695 300
rect 775 320 795 595
rect 775 25 795 300
rect 875 320 895 595
rect 875 25 895 300
rect 975 320 995 595
rect 1075 320 1095 595
rect 975 25 995 300
rect 1075 25 1095 300
rect 1175 320 1195 595
rect 1175 25 1195 300
rect 1275 320 1295 595
rect 1275 25 1295 300
rect 1375 320 1395 595
rect 1375 25 1395 300
rect 1475 320 1495 595
rect 1475 25 1495 300
rect 1575 320 1595 595
rect 1575 25 1595 300
<< pdiffc >>
rect -25 1055 -5 1330
rect -25 760 -5 1035
rect 75 1055 95 1330
rect 75 760 95 1035
rect 175 1055 195 1330
rect 175 760 195 1035
rect 275 1055 295 1330
rect 275 760 295 1035
rect 375 1055 395 1330
rect 375 760 395 1035
rect 475 1055 495 1330
rect 575 1055 595 1330
rect 475 760 495 1035
rect 575 760 595 1035
rect 675 1055 695 1330
rect 675 760 695 1035
rect 775 1055 795 1330
rect 775 760 795 1035
rect 875 1055 895 1330
rect 875 760 895 1035
rect 975 1055 995 1330
rect 975 760 995 1035
rect 1075 1055 1095 1330
rect 1075 760 1095 1035
rect 1175 1055 1195 1330
rect 1275 1055 1295 1330
rect 1175 760 1195 1035
rect 1275 760 1295 1035
rect 1375 1055 1395 1330
rect 1375 760 1395 1035
rect 1475 1055 1495 1330
rect 1475 760 1495 1035
rect 1575 1055 1595 1330
rect 1575 760 1595 1035
rect 1675 1055 1695 1330
rect 1675 760 1695 1035
rect 1775 1055 1795 1330
rect 1775 760 1795 1035
<< psubdiff >>
rect -90 595 -40 610
rect -90 320 -75 595
rect -55 320 -40 595
rect -90 300 -40 320
rect -90 25 -75 300
rect -55 25 -40 300
rect -90 10 -40 25
rect 510 595 560 610
rect 510 320 525 595
rect 545 320 560 595
rect 510 300 560 320
rect 510 25 525 300
rect 545 25 560 300
rect 510 10 560 25
rect 1010 595 1060 610
rect 1010 320 1025 595
rect 1045 320 1060 595
rect 1010 300 1060 320
rect 1010 25 1025 300
rect 1045 25 1060 300
rect 1010 10 1060 25
rect 1610 595 1660 610
rect 1610 320 1625 595
rect 1645 320 1660 595
rect 1610 300 1660 320
rect 1610 25 1625 300
rect 1645 25 1660 300
rect 1610 10 1660 25
<< nsubdiff >>
rect -90 1330 -40 1345
rect -90 1055 -75 1330
rect -55 1055 -40 1330
rect -90 1035 -40 1055
rect -90 760 -75 1035
rect -55 760 -40 1035
rect -90 745 -40 760
rect 510 1330 560 1345
rect 510 1055 525 1330
rect 545 1055 560 1330
rect 510 1035 560 1055
rect 510 760 525 1035
rect 545 760 560 1035
rect 510 745 560 760
rect 1210 1330 1260 1345
rect 1210 1055 1225 1330
rect 1245 1055 1260 1330
rect 1210 1035 1260 1055
rect 1210 760 1225 1035
rect 1245 760 1260 1035
rect 1210 745 1260 760
rect 1810 1330 1860 1345
rect 1810 1055 1825 1330
rect 1845 1055 1860 1330
rect 1810 1035 1860 1055
rect 1810 760 1825 1035
rect 1845 760 1860 1035
rect 1810 745 1860 760
<< psubdiffcont >>
rect -75 320 -55 595
rect -75 25 -55 300
rect 525 320 545 595
rect 525 25 545 300
rect 1025 320 1045 595
rect 1025 25 1045 300
rect 1625 320 1645 595
rect 1625 25 1645 300
<< nsubdiffcont >>
rect -75 1055 -55 1330
rect -75 760 -55 1035
rect 525 1055 545 1330
rect 525 760 545 1035
rect 1225 1055 1245 1330
rect 1225 760 1245 1035
rect 1825 1055 1845 1330
rect 1825 760 1845 1035
<< poly >>
rect 810 1385 1660 1400
rect 110 1360 760 1375
rect 10 1345 60 1360
rect 110 1345 160 1360
rect 210 1345 260 1360
rect 310 1345 360 1360
rect 410 1345 460 1360
rect 610 1345 660 1360
rect 710 1345 760 1360
rect 810 1345 860 1385
rect 910 1345 960 1360
rect 1010 1345 1060 1360
rect 1110 1345 1160 1385
rect 1310 1345 1360 1385
rect 1410 1345 1460 1360
rect 1510 1345 1560 1360
rect 1610 1345 1660 1385
rect 1710 1345 1760 1360
rect 10 730 60 745
rect 110 730 160 745
rect 210 730 260 745
rect 310 730 360 745
rect 410 730 460 745
rect 610 730 660 745
rect 710 730 760 745
rect 810 730 860 745
rect 910 730 960 745
rect 1010 730 1060 745
rect 1110 730 1160 745
rect 1310 730 1360 745
rect 1410 730 1460 745
rect 1510 730 1560 745
rect 1610 730 1660 745
rect 1710 730 1760 745
rect 910 705 1060 730
rect 1410 705 1560 730
rect 910 690 1560 705
rect 265 680 305 690
rect 265 665 275 680
rect 110 660 275 665
rect 295 665 305 680
rect 765 680 805 690
rect 765 665 775 680
rect 295 660 460 665
rect 110 650 460 660
rect 10 610 60 625
rect 110 610 160 650
rect 210 610 260 625
rect 310 610 360 625
rect 410 610 460 650
rect 610 660 775 665
rect 795 665 805 680
rect 795 660 1460 665
rect 610 650 1460 660
rect 610 610 660 650
rect 710 610 760 625
rect 810 610 860 625
rect 910 610 960 650
rect 1110 610 1160 650
rect 1210 610 1260 625
rect 1310 610 1360 625
rect 1410 610 1460 650
rect 1510 610 1560 625
rect 10 -5 60 10
rect 110 -5 160 10
rect -35 -15 60 -5
rect -35 -35 -25 -15
rect -5 -35 60 -15
rect -35 -45 60 -35
rect 210 -30 260 10
rect 310 -30 360 10
rect 410 -5 460 10
rect 610 -5 660 10
rect 710 -30 760 10
rect 810 -30 860 10
rect 910 -5 960 10
rect 1110 -5 1160 10
rect 1210 -30 1260 10
rect 1310 -30 1360 10
rect 1410 -5 1460 10
rect 1510 -5 1560 10
rect 210 -45 1360 -30
rect 1510 -15 1605 -5
rect 1510 -35 1575 -15
rect 1595 -35 1605 -15
rect 1510 -45 1605 -35
<< polycont >>
rect 275 660 295 680
rect 775 660 795 680
rect -25 -35 -5 -15
rect 1575 -35 1595 -15
<< locali >>
rect 685 1360 985 1380
rect 685 1340 705 1360
rect 965 1340 985 1360
rect -85 1330 5 1340
rect -85 1055 -75 1330
rect -55 1055 -25 1330
rect -5 1055 5 1330
rect -85 1035 5 1055
rect -85 760 -75 1035
rect -55 760 -25 1035
rect -5 760 5 1035
rect -85 750 5 760
rect 65 1330 105 1340
rect 65 1055 75 1330
rect 95 1055 105 1330
rect 65 1035 105 1055
rect 65 760 75 1035
rect 95 760 105 1035
rect 65 750 105 760
rect 165 1330 205 1340
rect 165 1055 175 1330
rect 195 1055 205 1330
rect 165 1035 205 1055
rect 165 760 175 1035
rect 195 760 205 1035
rect 165 750 205 760
rect 265 1330 305 1340
rect 265 1055 275 1330
rect 295 1055 305 1330
rect 265 1035 305 1055
rect 265 760 275 1035
rect 295 760 305 1035
rect 265 750 305 760
rect 365 1330 405 1340
rect 365 1055 375 1330
rect 395 1055 405 1330
rect 365 1035 405 1055
rect 365 760 375 1035
rect 395 760 405 1035
rect 365 750 405 760
rect 465 1330 605 1340
rect 465 1055 475 1330
rect 495 1055 525 1330
rect 545 1055 575 1330
rect 595 1055 605 1330
rect 465 1035 605 1055
rect 465 760 475 1035
rect 495 760 525 1035
rect 545 760 575 1035
rect 595 760 605 1035
rect 465 750 605 760
rect 665 1330 705 1340
rect 665 1055 675 1330
rect 695 1055 705 1330
rect 665 1035 705 1055
rect 665 760 675 1035
rect 695 760 705 1035
rect 665 750 705 760
rect 765 1330 805 1340
rect 765 1055 775 1330
rect 795 1055 805 1330
rect 765 1035 805 1055
rect 765 760 775 1035
rect 795 760 805 1035
rect 765 750 805 760
rect 865 1330 905 1340
rect 865 1055 875 1330
rect 895 1055 905 1330
rect 865 1035 905 1055
rect 865 760 875 1035
rect 895 760 905 1035
rect 865 750 905 760
rect 965 1330 1005 1340
rect 965 1055 975 1330
rect 995 1055 1005 1330
rect 965 1035 1005 1055
rect 965 760 975 1035
rect 995 760 1005 1035
rect 965 750 1005 760
rect 1065 1330 1105 1340
rect 1065 1055 1075 1330
rect 1095 1055 1105 1330
rect 1065 1035 1105 1055
rect 1065 760 1075 1035
rect 1095 760 1105 1035
rect 1065 750 1105 760
rect 1165 1330 1305 1340
rect 1165 1055 1175 1330
rect 1195 1055 1225 1330
rect 1245 1055 1275 1330
rect 1295 1055 1305 1330
rect 1165 1035 1305 1055
rect 1165 760 1175 1035
rect 1195 760 1225 1035
rect 1245 760 1275 1035
rect 1295 760 1305 1035
rect 1165 750 1305 760
rect 1365 1330 1405 1340
rect 1365 1055 1375 1330
rect 1395 1055 1405 1330
rect 1365 1035 1405 1055
rect 1365 760 1375 1035
rect 1395 760 1405 1035
rect 1365 750 1405 760
rect 1465 1330 1505 1340
rect 1465 1055 1475 1330
rect 1495 1055 1505 1330
rect 1465 1035 1505 1055
rect 1465 760 1475 1035
rect 1495 760 1505 1035
rect 1465 750 1505 760
rect 1565 1330 1605 1340
rect 1565 1055 1575 1330
rect 1595 1055 1605 1330
rect 1565 1035 1605 1055
rect 1565 760 1575 1035
rect 1595 760 1605 1035
rect 1565 750 1605 760
rect 1665 1330 1705 1340
rect 1665 1055 1675 1330
rect 1695 1055 1705 1330
rect 1665 1035 1705 1055
rect 1665 760 1675 1035
rect 1695 760 1705 1035
rect 1665 750 1705 760
rect 1765 1330 1855 1340
rect 1765 1055 1775 1330
rect 1795 1055 1825 1330
rect 1845 1055 1855 1330
rect 1765 1035 1855 1055
rect 1765 760 1775 1035
rect 1795 760 1825 1035
rect 1845 760 1855 1035
rect 1765 750 1855 760
rect 165 690 185 750
rect 365 690 385 750
rect 165 680 305 690
rect 165 670 275 680
rect 265 660 275 670
rect 295 660 305 680
rect 365 680 805 690
rect 365 670 775 680
rect 265 650 305 660
rect 765 660 775 670
rect 795 660 805 680
rect 765 650 805 660
rect 975 655 995 750
rect 275 605 295 650
rect 775 605 795 650
rect 975 635 1285 655
rect 1265 605 1285 635
rect -85 595 5 605
rect -85 320 -75 595
rect -55 320 -25 595
rect -5 320 5 595
rect -85 300 5 320
rect -85 25 -75 300
rect -55 25 -25 300
rect -5 25 5 300
rect -85 15 5 25
rect 65 595 105 605
rect 65 320 75 595
rect 95 320 105 595
rect 65 300 105 320
rect 65 25 75 300
rect 95 25 105 300
rect 65 15 105 25
rect 165 595 205 605
rect 165 320 175 595
rect 195 320 205 595
rect 165 300 205 320
rect 165 25 175 300
rect 195 25 205 300
rect 165 15 205 25
rect 265 595 305 605
rect 265 320 275 595
rect 295 320 305 595
rect 265 300 305 320
rect 265 25 275 300
rect 295 25 305 300
rect 265 15 305 25
rect 365 595 405 605
rect 365 320 375 595
rect 395 320 405 595
rect 365 300 405 320
rect 365 25 375 300
rect 395 25 405 300
rect 365 15 405 25
rect 465 595 605 605
rect 465 320 475 595
rect 495 320 525 595
rect 545 320 575 595
rect 595 320 605 595
rect 465 300 605 320
rect 465 25 475 300
rect 495 25 525 300
rect 545 25 575 300
rect 595 25 605 300
rect 465 15 605 25
rect 665 595 705 605
rect 665 320 675 595
rect 695 320 705 595
rect 665 300 705 320
rect 665 25 675 300
rect 695 25 705 300
rect 665 15 705 25
rect 765 595 805 605
rect 765 320 775 595
rect 795 320 805 595
rect 765 300 805 320
rect 765 25 775 300
rect 795 25 805 300
rect 765 15 805 25
rect 865 595 905 605
rect 865 320 875 595
rect 895 320 905 595
rect 865 300 905 320
rect 865 25 875 300
rect 895 25 905 300
rect 865 15 905 25
rect 965 595 1105 605
rect 965 320 975 595
rect 995 320 1025 595
rect 1045 320 1075 595
rect 1095 320 1105 595
rect 965 300 1105 320
rect 965 25 975 300
rect 995 25 1025 300
rect 1045 25 1075 300
rect 1095 25 1105 300
rect 965 15 1105 25
rect 1165 595 1205 605
rect 1165 320 1175 595
rect 1195 320 1205 595
rect 1165 300 1205 320
rect 1165 25 1175 300
rect 1195 25 1205 300
rect 1165 15 1205 25
rect 1265 595 1305 605
rect 1265 320 1275 595
rect 1295 320 1305 595
rect 1265 300 1305 320
rect 1265 25 1275 300
rect 1295 25 1305 300
rect 1265 15 1305 25
rect 1365 595 1405 605
rect 1365 320 1375 595
rect 1395 320 1405 595
rect 1365 300 1405 320
rect 1365 25 1375 300
rect 1395 25 1405 300
rect 1365 15 1405 25
rect 1465 595 1505 605
rect 1465 320 1475 595
rect 1495 320 1505 595
rect 1465 300 1505 320
rect 1465 25 1475 300
rect 1495 25 1505 300
rect 1465 15 1505 25
rect 1565 595 1655 605
rect 1565 320 1575 595
rect 1595 320 1625 595
rect 1645 320 1655 595
rect 1565 300 1655 320
rect 1565 25 1575 300
rect 1595 25 1625 300
rect 1645 25 1655 300
rect 1565 15 1655 25
rect -25 -5 -5 15
rect 185 -5 205 15
rect 365 -5 385 15
rect -35 -15 5 -5
rect -35 -35 -25 -15
rect -5 -35 5 -15
rect 185 -25 385 -5
rect 665 -5 685 15
rect 865 -5 885 15
rect 1575 -5 1595 15
rect 665 -25 885 -5
rect 1565 -15 1605 -5
rect -35 -45 5 -35
rect 1565 -35 1575 -15
rect 1595 -35 1605 -15
rect 1565 -45 1605 -35
<< end >>

magic
tech sky130A
timestamp 1699932530
<< nwell >>
rect -110 690 1880 1400
<< nmos >>
rect 10 -15 60 585
rect 110 -15 160 585
rect 210 -15 260 585
rect 310 -15 360 585
rect 410 -15 460 585
rect 610 -15 660 585
rect 710 -15 760 585
rect 810 -15 860 585
rect 910 -15 960 585
rect 1110 -15 1160 585
rect 1210 -15 1260 585
rect 1310 -15 1360 585
rect 1410 -15 1460 585
rect 1510 -15 1560 585
<< pmos >>
rect 10 745 60 1345
rect 110 745 160 1345
rect 210 745 260 1345
rect 310 745 360 1345
rect 410 745 460 1345
rect 610 745 660 1345
rect 710 745 760 1345
rect 810 745 860 1345
rect 910 745 960 1345
rect 1010 745 1060 1345
rect 1110 745 1160 1345
rect 1310 745 1360 1345
rect 1410 745 1460 1345
rect 1510 745 1560 1345
rect 1610 745 1660 1345
rect 1710 745 1760 1345
<< ndiff >>
rect -40 570 10 585
rect -40 295 -25 570
rect -5 295 10 570
rect -40 275 10 295
rect -40 0 -25 275
rect -5 0 10 275
rect -40 -15 10 0
rect 60 570 110 585
rect 60 295 75 570
rect 95 295 110 570
rect 60 275 110 295
rect 60 0 75 275
rect 95 0 110 275
rect 60 -15 110 0
rect 160 570 210 585
rect 160 295 175 570
rect 195 295 210 570
rect 160 275 210 295
rect 160 0 175 275
rect 195 0 210 275
rect 160 -15 210 0
rect 260 570 310 585
rect 260 295 275 570
rect 295 295 310 570
rect 260 275 310 295
rect 260 0 275 275
rect 295 0 310 275
rect 260 -15 310 0
rect 360 570 410 585
rect 360 295 375 570
rect 395 295 410 570
rect 360 275 410 295
rect 360 0 375 275
rect 395 0 410 275
rect 360 -15 410 0
rect 460 570 510 585
rect 560 570 610 585
rect 460 295 475 570
rect 495 295 510 570
rect 560 295 575 570
rect 595 295 610 570
rect 460 275 510 295
rect 560 275 610 295
rect 460 0 475 275
rect 495 0 510 275
rect 560 0 575 275
rect 595 0 610 275
rect 460 -15 510 0
rect 560 -15 610 0
rect 660 570 710 585
rect 660 295 675 570
rect 695 295 710 570
rect 660 275 710 295
rect 660 0 675 275
rect 695 0 710 275
rect 660 -15 710 0
rect 760 570 810 585
rect 760 295 775 570
rect 795 295 810 570
rect 760 275 810 295
rect 760 0 775 275
rect 795 0 810 275
rect 760 -15 810 0
rect 860 570 910 585
rect 860 295 875 570
rect 895 295 910 570
rect 860 275 910 295
rect 860 0 875 275
rect 895 0 910 275
rect 860 -15 910 0
rect 960 570 1010 585
rect 1060 570 1110 585
rect 960 295 975 570
rect 995 295 1010 570
rect 1060 295 1075 570
rect 1095 295 1110 570
rect 960 275 1010 295
rect 1060 275 1110 295
rect 960 0 975 275
rect 995 0 1010 275
rect 1060 0 1075 275
rect 1095 0 1110 275
rect 960 -15 1010 0
rect 1060 -15 1110 0
rect 1160 570 1210 585
rect 1160 295 1175 570
rect 1195 295 1210 570
rect 1160 275 1210 295
rect 1160 0 1175 275
rect 1195 0 1210 275
rect 1160 -15 1210 0
rect 1260 570 1310 585
rect 1260 295 1275 570
rect 1295 295 1310 570
rect 1260 275 1310 295
rect 1260 0 1275 275
rect 1295 0 1310 275
rect 1260 -15 1310 0
rect 1360 570 1410 585
rect 1360 295 1375 570
rect 1395 295 1410 570
rect 1360 275 1410 295
rect 1360 0 1375 275
rect 1395 0 1410 275
rect 1360 -15 1410 0
rect 1460 570 1510 585
rect 1460 295 1475 570
rect 1495 295 1510 570
rect 1460 275 1510 295
rect 1460 0 1475 275
rect 1495 0 1510 275
rect 1460 -15 1510 0
rect 1560 570 1610 585
rect 1560 295 1575 570
rect 1595 295 1610 570
rect 1560 275 1610 295
rect 1560 0 1575 275
rect 1595 0 1610 275
rect 1560 -15 1610 0
<< pdiff >>
rect -40 1330 10 1345
rect -40 1055 -25 1330
rect -5 1055 10 1330
rect -40 1035 10 1055
rect -40 760 -25 1035
rect -5 760 10 1035
rect -40 745 10 760
rect 60 1330 110 1345
rect 60 1055 75 1330
rect 95 1055 110 1330
rect 60 1035 110 1055
rect 60 760 75 1035
rect 95 760 110 1035
rect 60 745 110 760
rect 160 1330 210 1345
rect 160 1055 175 1330
rect 195 1055 210 1330
rect 160 1035 210 1055
rect 160 760 175 1035
rect 195 760 210 1035
rect 160 745 210 760
rect 260 1330 310 1345
rect 260 1055 275 1330
rect 295 1055 310 1330
rect 260 1035 310 1055
rect 260 760 275 1035
rect 295 760 310 1035
rect 260 745 310 760
rect 360 1330 410 1345
rect 360 1055 375 1330
rect 395 1055 410 1330
rect 360 1035 410 1055
rect 360 760 375 1035
rect 395 760 410 1035
rect 360 745 410 760
rect 460 1330 510 1345
rect 560 1330 610 1345
rect 460 1055 475 1330
rect 495 1055 510 1330
rect 560 1055 575 1330
rect 595 1055 610 1330
rect 460 1035 510 1055
rect 560 1035 610 1055
rect 460 760 475 1035
rect 495 760 510 1035
rect 560 760 575 1035
rect 595 760 610 1035
rect 460 745 510 760
rect 560 745 610 760
rect 660 1330 710 1345
rect 660 1055 675 1330
rect 695 1055 710 1330
rect 660 1035 710 1055
rect 660 760 675 1035
rect 695 760 710 1035
rect 660 745 710 760
rect 760 1330 810 1345
rect 760 1055 775 1330
rect 795 1055 810 1330
rect 760 1035 810 1055
rect 760 760 775 1035
rect 795 760 810 1035
rect 760 745 810 760
rect 860 1330 910 1345
rect 860 1055 875 1330
rect 895 1055 910 1330
rect 860 1035 910 1055
rect 860 760 875 1035
rect 895 760 910 1035
rect 860 745 910 760
rect 960 1330 1010 1345
rect 960 1055 975 1330
rect 995 1055 1010 1330
rect 960 1035 1010 1055
rect 960 760 975 1035
rect 995 760 1010 1035
rect 960 745 1010 760
rect 1060 1330 1110 1345
rect 1060 1055 1075 1330
rect 1095 1055 1110 1330
rect 1060 1035 1110 1055
rect 1060 760 1075 1035
rect 1095 760 1110 1035
rect 1060 745 1110 760
rect 1160 1330 1210 1345
rect 1260 1330 1310 1345
rect 1160 1055 1175 1330
rect 1195 1055 1210 1330
rect 1260 1055 1275 1330
rect 1295 1055 1310 1330
rect 1160 1035 1210 1055
rect 1260 1035 1310 1055
rect 1160 760 1175 1035
rect 1195 760 1210 1035
rect 1260 760 1275 1035
rect 1295 760 1310 1035
rect 1160 745 1210 760
rect 1260 745 1310 760
rect 1360 1330 1410 1345
rect 1360 1055 1375 1330
rect 1395 1055 1410 1330
rect 1360 1035 1410 1055
rect 1360 760 1375 1035
rect 1395 760 1410 1035
rect 1360 745 1410 760
rect 1460 1330 1510 1345
rect 1460 1055 1475 1330
rect 1495 1055 1510 1330
rect 1460 1035 1510 1055
rect 1460 760 1475 1035
rect 1495 760 1510 1035
rect 1460 745 1510 760
rect 1560 1330 1610 1345
rect 1560 1055 1575 1330
rect 1595 1055 1610 1330
rect 1560 1035 1610 1055
rect 1560 760 1575 1035
rect 1595 760 1610 1035
rect 1560 745 1610 760
rect 1660 1330 1710 1345
rect 1660 1055 1675 1330
rect 1695 1055 1710 1330
rect 1660 1035 1710 1055
rect 1660 760 1675 1035
rect 1695 760 1710 1035
rect 1660 745 1710 760
rect 1760 1330 1810 1345
rect 1760 1055 1775 1330
rect 1795 1055 1810 1330
rect 1760 1035 1810 1055
rect 1760 760 1775 1035
rect 1795 760 1810 1035
rect 1760 745 1810 760
<< ndiffc >>
rect -25 295 -5 570
rect -25 0 -5 275
rect 75 295 95 570
rect 75 0 95 275
rect 175 295 195 570
rect 175 0 195 275
rect 275 295 295 570
rect 275 0 295 275
rect 375 295 395 570
rect 375 0 395 275
rect 475 295 495 570
rect 575 295 595 570
rect 475 0 495 275
rect 575 0 595 275
rect 675 295 695 570
rect 675 0 695 275
rect 775 295 795 570
rect 775 0 795 275
rect 875 295 895 570
rect 875 0 895 275
rect 975 295 995 570
rect 1075 295 1095 570
rect 975 0 995 275
rect 1075 0 1095 275
rect 1175 295 1195 570
rect 1175 0 1195 275
rect 1275 295 1295 570
rect 1275 0 1295 275
rect 1375 295 1395 570
rect 1375 0 1395 275
rect 1475 295 1495 570
rect 1475 0 1495 275
rect 1575 295 1595 570
rect 1575 0 1595 275
<< pdiffc >>
rect -25 1055 -5 1330
rect -25 760 -5 1035
rect 75 1055 95 1330
rect 75 760 95 1035
rect 175 1055 195 1330
rect 175 760 195 1035
rect 275 1055 295 1330
rect 275 760 295 1035
rect 375 1055 395 1330
rect 375 760 395 1035
rect 475 1055 495 1330
rect 575 1055 595 1330
rect 475 760 495 1035
rect 575 760 595 1035
rect 675 1055 695 1330
rect 675 760 695 1035
rect 775 1055 795 1330
rect 775 760 795 1035
rect 875 1055 895 1330
rect 875 760 895 1035
rect 975 1055 995 1330
rect 975 760 995 1035
rect 1075 1055 1095 1330
rect 1075 760 1095 1035
rect 1175 1055 1195 1330
rect 1275 1055 1295 1330
rect 1175 760 1195 1035
rect 1275 760 1295 1035
rect 1375 1055 1395 1330
rect 1375 760 1395 1035
rect 1475 1055 1495 1330
rect 1475 760 1495 1035
rect 1575 1055 1595 1330
rect 1575 760 1595 1035
rect 1675 1055 1695 1330
rect 1675 760 1695 1035
rect 1775 1055 1795 1330
rect 1775 760 1795 1035
<< psubdiff >>
rect -90 570 -40 585
rect -90 295 -75 570
rect -55 295 -40 570
rect -90 275 -40 295
rect -90 0 -75 275
rect -55 0 -40 275
rect -90 -15 -40 0
rect 510 570 560 585
rect 510 295 525 570
rect 545 295 560 570
rect 510 275 560 295
rect 510 0 525 275
rect 545 0 560 275
rect 510 -15 560 0
rect 1010 570 1060 585
rect 1010 295 1025 570
rect 1045 295 1060 570
rect 1010 275 1060 295
rect 1010 0 1025 275
rect 1045 0 1060 275
rect 1010 -15 1060 0
rect 1610 570 1660 585
rect 1610 295 1625 570
rect 1645 295 1660 570
rect 1610 275 1660 295
rect 1610 0 1625 275
rect 1645 0 1660 275
rect 1610 -15 1660 0
<< nsubdiff >>
rect -90 1330 -40 1345
rect -90 1055 -75 1330
rect -55 1055 -40 1330
rect -90 1035 -40 1055
rect -90 760 -75 1035
rect -55 760 -40 1035
rect -90 745 -40 760
rect 510 1330 560 1345
rect 510 1055 525 1330
rect 545 1055 560 1330
rect 510 1035 560 1055
rect 510 760 525 1035
rect 545 760 560 1035
rect 510 745 560 760
rect 1210 1330 1260 1345
rect 1210 1055 1225 1330
rect 1245 1055 1260 1330
rect 1210 1035 1260 1055
rect 1210 760 1225 1035
rect 1245 760 1260 1035
rect 1210 745 1260 760
rect 1810 1330 1860 1345
rect 1810 1055 1825 1330
rect 1845 1055 1860 1330
rect 1810 1035 1860 1055
rect 1810 760 1825 1035
rect 1845 760 1860 1035
rect 1810 745 1860 760
<< psubdiffcont >>
rect -75 295 -55 570
rect -75 0 -55 275
rect 525 295 545 570
rect 525 0 545 275
rect 1025 295 1045 570
rect 1025 0 1045 275
rect 1625 295 1645 570
rect 1625 0 1645 275
<< nsubdiffcont >>
rect -75 1055 -55 1330
rect -75 760 -55 1035
rect 525 1055 545 1330
rect 525 760 545 1035
rect 1225 1055 1245 1330
rect 1225 760 1245 1035
rect 1825 1055 1845 1330
rect 1825 760 1845 1035
<< poly >>
rect -95 1425 125 1440
rect -95 1410 -80 1425
rect -140 1395 -80 1410
rect -35 1390 5 1400
rect -35 1370 -25 1390
rect -5 1380 5 1390
rect -5 1370 60 1380
rect -35 1360 60 1370
rect 10 1345 60 1360
rect 110 1375 125 1425
rect 810 1390 1660 1400
rect 110 1360 760 1375
rect 110 1345 160 1360
rect 210 1345 260 1360
rect 310 1345 360 1360
rect 410 1345 460 1360
rect 610 1345 660 1360
rect 710 1345 760 1360
rect 810 1370 825 1390
rect 845 1385 1660 1390
rect 845 1370 860 1385
rect 810 1345 860 1370
rect 910 1345 960 1360
rect 1010 1345 1060 1360
rect 1110 1345 1160 1385
rect 1310 1345 1360 1385
rect 1410 1345 1460 1360
rect 1510 1345 1560 1360
rect 1610 1345 1660 1385
rect 1765 1390 1805 1400
rect 1765 1375 1775 1390
rect 1745 1370 1775 1375
rect 1795 1370 1805 1390
rect 1745 1360 1805 1370
rect 1710 1345 1760 1360
rect 10 730 60 745
rect 110 730 160 745
rect 210 730 260 745
rect 310 730 360 745
rect 410 730 460 745
rect 610 730 660 745
rect 710 730 760 745
rect 810 730 860 745
rect 910 730 960 745
rect 1010 730 1060 745
rect 1110 730 1160 745
rect 1310 730 1360 745
rect 1410 730 1460 745
rect 1510 730 1560 745
rect 1610 730 1660 745
rect 1710 730 1760 745
rect 910 705 1060 730
rect 1410 705 1560 730
rect -140 690 1560 705
rect 265 655 305 665
rect 265 640 275 655
rect 110 635 275 640
rect 295 640 305 655
rect 765 655 805 665
rect 765 640 775 655
rect 295 635 460 640
rect 110 625 460 635
rect 10 585 60 600
rect 110 585 160 625
rect 210 585 260 600
rect 310 585 360 600
rect 410 585 460 625
rect 610 635 775 640
rect 795 640 805 655
rect 795 635 1460 640
rect 610 625 1460 635
rect 610 585 660 625
rect 710 585 760 600
rect 810 585 860 600
rect 910 585 960 625
rect 1110 585 1160 625
rect 1210 585 1260 600
rect 1310 585 1360 600
rect 1410 585 1460 625
rect 1510 585 1560 600
rect 10 -30 60 -15
rect 110 -30 160 -15
rect -35 -40 60 -30
rect -35 -60 -25 -40
rect -5 -60 60 -40
rect -35 -70 60 -60
rect 210 -55 260 -15
rect 310 -55 360 -15
rect 410 -30 460 -15
rect 610 -30 660 -15
rect 710 -55 760 -15
rect 810 -55 860 -15
rect 910 -30 960 -15
rect 1110 -30 1160 -15
rect 1210 -55 1260 -15
rect 1310 -55 1360 -15
rect 1410 -30 1460 -15
rect 1510 -30 1560 -15
rect 210 -70 1360 -55
rect 1510 -40 1605 -30
rect 1510 -60 1575 -40
rect 1595 -60 1605 -40
rect 1510 -70 1605 -60
rect 210 -115 225 -70
rect -140 -130 225 -115
<< polycont >>
rect -25 1370 -5 1390
rect 825 1370 845 1390
rect 1775 1370 1795 1390
rect 275 635 295 655
rect 775 635 795 655
rect -25 -60 -5 -40
rect 1575 -60 1595 -40
<< locali >>
rect -140 1420 1485 1440
rect -35 1390 5 1400
rect -35 1370 -25 1390
rect -5 1370 5 1390
rect 815 1390 855 1400
rect 815 1380 825 1390
rect -35 1360 5 1370
rect 685 1370 825 1380
rect 845 1380 855 1390
rect 845 1370 985 1380
rect 685 1360 985 1370
rect -25 1340 -5 1360
rect 685 1340 705 1360
rect 965 1340 985 1360
rect 1465 1340 1485 1420
rect 1765 1390 1805 1400
rect 1765 1370 1775 1390
rect 1795 1370 1805 1390
rect 1765 1360 1805 1370
rect 1775 1340 1795 1360
rect -85 1330 5 1340
rect -85 1055 -75 1330
rect -55 1055 -25 1330
rect -5 1055 5 1330
rect -85 1035 5 1055
rect -85 760 -75 1035
rect -55 760 -25 1035
rect -5 760 5 1035
rect -85 750 5 760
rect 65 1330 105 1340
rect 65 1055 75 1330
rect 95 1055 105 1330
rect 65 1035 105 1055
rect 65 760 75 1035
rect 95 760 105 1035
rect 65 750 105 760
rect 165 1330 205 1340
rect 165 1055 175 1330
rect 195 1055 205 1330
rect 165 1035 205 1055
rect 165 760 175 1035
rect 195 760 205 1035
rect 165 750 205 760
rect 265 1330 305 1340
rect 265 1055 275 1330
rect 295 1055 305 1330
rect 265 1035 305 1055
rect 265 760 275 1035
rect 295 760 305 1035
rect 265 750 305 760
rect 365 1330 405 1340
rect 365 1055 375 1330
rect 395 1055 405 1330
rect 365 1035 405 1055
rect 365 760 375 1035
rect 395 760 405 1035
rect 365 750 405 760
rect 465 1330 605 1340
rect 465 1055 475 1330
rect 495 1055 525 1330
rect 545 1055 575 1330
rect 595 1055 605 1330
rect 465 1035 605 1055
rect 465 760 475 1035
rect 495 760 525 1035
rect 545 760 575 1035
rect 595 760 605 1035
rect 465 750 605 760
rect 665 1330 705 1340
rect 665 1055 675 1330
rect 695 1055 705 1330
rect 665 1035 705 1055
rect 665 760 675 1035
rect 695 760 705 1035
rect 665 750 705 760
rect 765 1330 805 1340
rect 765 1055 775 1330
rect 795 1055 805 1330
rect 765 1035 805 1055
rect 765 760 775 1035
rect 795 760 805 1035
rect 765 750 805 760
rect 865 1330 905 1340
rect 865 1055 875 1330
rect 895 1055 905 1330
rect 865 1035 905 1055
rect 865 760 875 1035
rect 895 760 905 1035
rect 865 750 905 760
rect 965 1330 1005 1340
rect 965 1055 975 1330
rect 995 1055 1005 1330
rect 965 1035 1005 1055
rect 965 760 975 1035
rect 995 760 1005 1035
rect 965 750 1005 760
rect 1065 1330 1105 1340
rect 1065 1055 1075 1330
rect 1095 1055 1105 1330
rect 1065 1035 1105 1055
rect 1065 760 1075 1035
rect 1095 760 1105 1035
rect 1065 750 1105 760
rect 1165 1330 1305 1340
rect 1165 1055 1175 1330
rect 1195 1055 1225 1330
rect 1245 1055 1275 1330
rect 1295 1055 1305 1330
rect 1165 1035 1305 1055
rect 1165 760 1175 1035
rect 1195 760 1225 1035
rect 1245 760 1275 1035
rect 1295 760 1305 1035
rect 1165 750 1305 760
rect 1365 1330 1405 1340
rect 1365 1055 1375 1330
rect 1395 1055 1405 1330
rect 1365 1035 1405 1055
rect 1365 760 1375 1035
rect 1395 760 1405 1035
rect 1365 750 1405 760
rect 1465 1330 1505 1340
rect 1465 1055 1475 1330
rect 1495 1055 1505 1330
rect 1465 1035 1505 1055
rect 1465 760 1475 1035
rect 1495 760 1505 1035
rect 1465 750 1505 760
rect 1565 1330 1605 1340
rect 1565 1055 1575 1330
rect 1595 1055 1605 1330
rect 1565 1035 1605 1055
rect 1565 760 1575 1035
rect 1595 760 1605 1035
rect 1565 750 1605 760
rect 1665 1330 1705 1340
rect 1665 1055 1675 1330
rect 1695 1055 1705 1330
rect 1665 1035 1705 1055
rect 1665 760 1675 1035
rect 1695 760 1705 1035
rect 1665 750 1705 760
rect 1765 1330 1855 1340
rect 1765 1055 1775 1330
rect 1795 1055 1825 1330
rect 1845 1055 1855 1330
rect 1765 1035 1855 1055
rect 1765 760 1775 1035
rect 1795 760 1825 1035
rect 1845 760 1855 1035
rect 1765 750 1855 760
rect 165 665 185 750
rect 365 665 385 750
rect 165 655 305 665
rect 165 645 275 655
rect 265 635 275 645
rect 295 635 305 655
rect 365 655 805 665
rect 365 645 775 655
rect 265 625 305 635
rect 765 635 775 645
rect 795 635 805 655
rect 765 625 805 635
rect 975 630 995 750
rect 275 580 295 625
rect 775 580 795 625
rect 975 610 1880 630
rect 1265 580 1285 610
rect -85 570 5 580
rect -85 295 -75 570
rect -55 295 -25 570
rect -5 295 5 570
rect -85 275 5 295
rect -85 0 -75 275
rect -55 0 -25 275
rect -5 0 5 275
rect -85 -10 5 0
rect 65 570 105 580
rect 65 295 75 570
rect 95 295 105 570
rect 65 275 105 295
rect 65 0 75 275
rect 95 0 105 275
rect 65 -10 105 0
rect 165 570 205 580
rect 165 295 175 570
rect 195 295 205 570
rect 165 275 205 295
rect 165 0 175 275
rect 195 0 205 275
rect 165 -10 205 0
rect 265 570 305 580
rect 265 295 275 570
rect 295 295 305 570
rect 265 275 305 295
rect 265 0 275 275
rect 295 0 305 275
rect 265 -10 305 0
rect 365 570 405 580
rect 365 295 375 570
rect 395 295 405 570
rect 365 275 405 295
rect 365 0 375 275
rect 395 0 405 275
rect 365 -10 405 0
rect 465 570 605 580
rect 465 295 475 570
rect 495 295 525 570
rect 545 295 575 570
rect 595 295 605 570
rect 465 275 605 295
rect 465 0 475 275
rect 495 0 525 275
rect 545 0 575 275
rect 595 0 605 275
rect 465 -10 605 0
rect 665 570 705 580
rect 665 295 675 570
rect 695 295 705 570
rect 665 275 705 295
rect 665 0 675 275
rect 695 0 705 275
rect 665 -10 705 0
rect 765 570 805 580
rect 765 295 775 570
rect 795 295 805 570
rect 765 275 805 295
rect 765 0 775 275
rect 795 0 805 275
rect 765 -10 805 0
rect 865 570 905 580
rect 865 295 875 570
rect 895 295 905 570
rect 865 275 905 295
rect 865 0 875 275
rect 895 0 905 275
rect 865 -10 905 0
rect 965 570 1105 580
rect 965 295 975 570
rect 995 295 1025 570
rect 1045 295 1075 570
rect 1095 295 1105 570
rect 965 275 1105 295
rect 965 0 975 275
rect 995 0 1025 275
rect 1045 0 1075 275
rect 1095 0 1105 275
rect 965 -10 1105 0
rect 1165 570 1205 580
rect 1165 295 1175 570
rect 1195 295 1205 570
rect 1165 275 1205 295
rect 1165 0 1175 275
rect 1195 0 1205 275
rect 1165 -10 1205 0
rect 1265 570 1305 580
rect 1265 295 1275 570
rect 1295 295 1305 570
rect 1265 275 1305 295
rect 1265 0 1275 275
rect 1295 0 1305 275
rect 1265 -10 1305 0
rect 1365 570 1405 580
rect 1365 295 1375 570
rect 1395 295 1405 570
rect 1365 275 1405 295
rect 1365 0 1375 275
rect 1395 0 1405 275
rect 1365 -10 1405 0
rect 1465 570 1505 580
rect 1465 295 1475 570
rect 1495 295 1505 570
rect 1465 275 1505 295
rect 1465 0 1475 275
rect 1495 0 1505 275
rect 1465 -10 1505 0
rect 1565 570 1655 580
rect 1565 295 1575 570
rect 1595 295 1625 570
rect 1645 295 1655 570
rect 1565 275 1655 295
rect 1565 0 1575 275
rect 1595 0 1625 275
rect 1645 0 1655 275
rect 1565 -10 1655 0
rect -25 -30 -5 -10
rect 185 -30 205 -10
rect 365 -30 385 -10
rect -35 -40 5 -30
rect -35 -60 -25 -40
rect -5 -60 5 -40
rect -35 -70 5 -60
rect 185 -50 385 -30
rect 665 -30 685 -10
rect 865 -30 885 -10
rect 1575 -30 1595 -10
rect 665 -50 885 -30
rect 1565 -40 1605 -30
rect 185 -90 205 -50
rect -140 -110 205 -90
rect 665 -130 685 -50
rect 1565 -60 1575 -40
rect 1595 -60 1605 -40
rect 1565 -70 1605 -60
rect -140 -150 685 -130
<< viali >>
rect -75 1055 -55 1330
rect -25 1055 -5 1330
rect -75 760 -55 1035
rect -25 760 -5 1035
rect 75 1055 95 1330
rect 75 760 95 1035
rect 275 1055 295 1330
rect 275 760 295 1035
rect 475 1055 495 1330
rect 525 1055 545 1330
rect 575 1055 595 1330
rect 475 760 495 1035
rect 525 760 545 1035
rect 575 760 595 1035
rect 775 1055 795 1330
rect 775 760 795 1035
rect 1175 1055 1195 1330
rect 1225 1055 1245 1330
rect 1275 1055 1295 1330
rect 1175 760 1195 1035
rect 1225 760 1245 1035
rect 1275 760 1295 1035
rect 1675 1055 1695 1330
rect 1675 760 1695 1035
rect 1775 1055 1795 1330
rect 1825 1055 1845 1330
rect 1775 760 1795 1035
rect 1825 760 1845 1035
rect -75 295 -55 570
rect -25 295 -5 570
rect -75 0 -55 275
rect -25 0 -5 275
rect 75 295 95 570
rect 75 0 95 275
rect 475 295 495 570
rect 525 295 545 570
rect 575 295 595 570
rect 475 0 495 275
rect 525 0 545 275
rect 575 0 595 275
rect 975 295 995 570
rect 1025 295 1045 570
rect 1075 295 1095 570
rect 975 0 995 275
rect 1025 0 1045 275
rect 1075 0 1095 275
rect 1475 295 1495 570
rect 1475 0 1495 275
rect 1575 295 1595 570
rect 1625 295 1645 570
rect 1575 0 1595 275
rect 1625 0 1645 275
<< metal1 >>
rect -140 1330 1860 1340
rect -140 1055 -75 1330
rect -55 1055 -25 1330
rect -5 1055 75 1330
rect 95 1055 275 1330
rect 295 1055 475 1330
rect 495 1055 525 1330
rect 545 1055 575 1330
rect 595 1055 775 1330
rect 795 1055 1175 1330
rect 1195 1055 1225 1330
rect 1245 1055 1275 1330
rect 1295 1055 1675 1330
rect 1695 1055 1775 1330
rect 1795 1055 1825 1330
rect 1845 1055 1860 1330
rect -140 1035 1860 1055
rect -140 760 -75 1035
rect -55 760 -25 1035
rect -5 760 75 1035
rect 95 760 275 1035
rect 295 760 475 1035
rect 495 760 525 1035
rect 545 760 575 1035
rect 595 760 775 1035
rect 795 760 1175 1035
rect 1195 760 1225 1035
rect 1245 760 1275 1035
rect 1295 760 1675 1035
rect 1695 760 1775 1035
rect 1795 760 1825 1035
rect 1845 760 1860 1035
rect -140 750 1860 760
rect -140 570 1660 580
rect -140 295 -75 570
rect -55 295 -25 570
rect -5 295 75 570
rect 95 295 475 570
rect 495 295 525 570
rect 545 295 575 570
rect 595 295 975 570
rect 995 295 1025 570
rect 1045 295 1075 570
rect 1095 295 1475 570
rect 1495 295 1575 570
rect 1595 295 1625 570
rect 1645 295 1660 570
rect -140 275 1660 295
rect -140 0 -75 275
rect -55 0 -25 275
rect -5 0 75 275
rect 95 0 475 275
rect 495 0 525 275
rect 545 0 575 275
rect 595 0 975 275
rect 995 0 1025 275
rect 1045 0 1075 275
rect 1095 0 1475 275
rect 1495 0 1575 275
rect 1595 0 1625 275
rect 1645 0 1660 275
rect -140 -10 1660 0
<< labels >>
flabel locali -140 1430 -140 1430 7 FreeSans 160 0 0 0 Vbias
port 1 w
flabel metal1 -140 1045 -140 1045 7 FreeSans 160 0 0 0 VDD
port 2 w
flabel poly -140 1400 -140 1400 7 FreeSans 160 0 0 0 Vbp
port 7 w
flabel locali 1880 620 1880 620 3 FreeSans 160 0 0 0 Iout
port 6 e
flabel locali -140 -140 -140 -140 7 FreeSans 160 0 0 0 Idac
port 5 w
flabel locali -140 -100 -140 -100 7 FreeSans 160 0 0 0 Idump
port 4 w
flabel metal1 -140 285 -140 285 7 FreeSans 160 0 0 0 GND
port 3 w
flabel poly -140 695 -140 695 7 FreeSans 160 0 0 0 Vcp
port 8 w
flabel poly -140 -125 -140 -125 7 FreeSans 160 0 0 0 Vbn
port 9 w
<< end >>
